parameter CFIFO_DEPTH = 256;
