library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity rom16k is
    Port ( CLK : in  STD_LOGIC;
             A : in  STD_LOGIC_VECTOR (13 downto 0);
		   DIN : in  STD_LOGIC_VECTOR (7 downto 0);
          DOUT : out STD_LOGIC_VECTOR (7 downto 0);
			WR : in  STD_LOGIC);
				
end rom16k;

architecture Behavioral of rom16k is

type
  romarray is array(0 to 16383) of std_logic_vector(7 downto 0);

signal myROM : romarray := (

x"F3",x"AF",x"11",x"FF",x"FF",x"C3",x"8E",x"38",x"2A",x"5D",x"5C",x"22",x"5F",x"5C",x"18",x"43",
x"C3",x"F2",x"15",x"FF",x"FF",x"FF",x"FF",x"FF",x"2A",x"5D",x"5C",x"7E",x"CD",x"7D",x"00",x"D0",
x"CD",x"74",x"00",x"18",x"F7",x"FF",x"FF",x"FF",x"C3",x"5B",x"33",x"FF",x"FF",x"FF",x"FF",x"FF",
x"C5",x"2A",x"61",x"5C",x"E5",x"C3",x"9E",x"16",x"F5",x"E5",x"2A",x"78",x"5C",x"23",x"22",x"78",
x"5C",x"7C",x"B5",x"20",x"03",x"FD",x"34",x"40",x"C5",x"D5",x"CD",x"BF",x"02",x"D1",x"C1",x"E1",
x"F1",x"FB",x"C9",x"E1",x"6E",x"FD",x"75",x"00",x"ED",x"7B",x"3D",x"5C",x"C3",x"C5",x"16",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"F5",x"E5",x"2A",x"B0",x"5C",x"7C",x"B5",x"20",x"01",x"E9",
x"E1",x"F1",x"ED",x"45",x"2A",x"5D",x"5C",x"23",x"22",x"5D",x"5C",x"7E",x"C9",x"FE",x"21",x"D0",
x"FE",x"0D",x"C8",x"FE",x"10",x"D8",x"FE",x"18",x"3F",x"D8",x"23",x"FE",x"16",x"38",x"01",x"23",
x"37",x"22",x"5D",x"5C",x"C9",x"BF",x"52",x"4E",x"C4",x"49",x"4E",x"4B",x"45",x"59",x"A4",x"50",
x"C9",x"46",x"CE",x"50",x"4F",x"49",x"4E",x"D4",x"53",x"43",x"52",x"45",x"45",x"4E",x"A4",x"41",
x"54",x"54",x"D2",x"41",x"D4",x"54",x"41",x"C2",x"56",x"41",x"4C",x"A4",x"43",x"4F",x"44",x"C5",
x"56",x"41",x"CC",x"4C",x"45",x"CE",x"53",x"49",x"CE",x"43",x"4F",x"D3",x"54",x"41",x"CE",x"41",
x"53",x"CE",x"41",x"43",x"D3",x"41",x"54",x"CE",x"4C",x"CE",x"45",x"58",x"D0",x"49",x"4E",x"D4",
x"53",x"51",x"D2",x"53",x"47",x"CE",x"41",x"42",x"D3",x"50",x"45",x"45",x"CB",x"49",x"CE",x"55",
x"53",x"D2",x"53",x"54",x"52",x"A4",x"43",x"48",x"52",x"A4",x"4E",x"4F",x"D4",x"42",x"49",x"CE",
x"4F",x"D2",x"41",x"4E",x"C4",x"3C",x"BD",x"3E",x"BD",x"3C",x"BE",x"4C",x"49",x"4E",x"C5",x"54",
x"48",x"45",x"CE",x"54",x"CF",x"53",x"54",x"45",x"D0",x"44",x"45",x"46",x"20",x"46",x"CE",x"43",
x"41",x"D4",x"46",x"4F",x"52",x"4D",x"41",x"D4",x"4D",x"4F",x"56",x"C5",x"45",x"52",x"41",x"53",
x"C5",x"4F",x"50",x"45",x"4E",x"20",x"A3",x"43",x"4C",x"4F",x"53",x"45",x"20",x"A3",x"4D",x"45",
x"52",x"47",x"C5",x"56",x"45",x"52",x"49",x"46",x"D9",x"42",x"45",x"45",x"D0",x"43",x"49",x"52",
x"43",x"4C",x"C5",x"49",x"4E",x"CB",x"50",x"41",x"50",x"45",x"D2",x"46",x"4C",x"41",x"53",x"C8",
x"42",x"52",x"49",x"47",x"48",x"D4",x"49",x"4E",x"56",x"45",x"52",x"53",x"C5",x"4F",x"56",x"45",
x"D2",x"4F",x"55",x"D4",x"4C",x"50",x"52",x"49",x"4E",x"D4",x"4C",x"4C",x"49",x"53",x"D4",x"53",
x"54",x"4F",x"D0",x"52",x"45",x"41",x"C4",x"44",x"41",x"54",x"C1",x"52",x"45",x"53",x"54",x"4F",
x"52",x"C5",x"4E",x"45",x"D7",x"42",x"4F",x"52",x"44",x"45",x"D2",x"43",x"4F",x"4E",x"54",x"49",
x"4E",x"55",x"C5",x"44",x"49",x"CD",x"52",x"45",x"CD",x"46",x"4F",x"D2",x"47",x"4F",x"20",x"54",
x"CF",x"47",x"4F",x"20",x"53",x"55",x"C2",x"49",x"4E",x"50",x"55",x"D4",x"4C",x"4F",x"41",x"C4",
x"4C",x"49",x"53",x"D4",x"4C",x"45",x"D4",x"50",x"41",x"55",x"53",x"C5",x"4E",x"45",x"58",x"D4",
x"50",x"4F",x"4B",x"C5",x"50",x"52",x"49",x"4E",x"D4",x"50",x"4C",x"4F",x"D4",x"52",x"55",x"CE",
x"53",x"41",x"56",x"C5",x"52",x"41",x"4E",x"44",x"4F",x"4D",x"49",x"5A",x"C5",x"49",x"C6",x"43",
x"4C",x"D3",x"44",x"52",x"41",x"D7",x"43",x"4C",x"45",x"41",x"D2",x"52",x"45",x"54",x"55",x"52",
x"CE",x"43",x"4D",x"C4",x"D9",x"42",x"48",x"59",x"36",x"35",x"54",x"47",x"56",x"4E",x"4A",x"55",
x"37",x"34",x"52",x"46",x"43",x"4D",x"4B",x"49",x"38",x"33",x"45",x"44",x"58",x"0E",x"4C",x"4F",
x"39",x"32",x"57",x"53",x"5A",x"20",x"0D",x"50",x"30",x"31",x"51",x"41",x"E3",x"C4",x"E0",x"E4",
x"B4",x"BC",x"BD",x"BB",x"AF",x"B0",x"B1",x"C0",x"A7",x"A6",x"BE",x"AD",x"B2",x"BA",x"E5",x"A5",
x"C2",x"E1",x"B3",x"B9",x"C1",x"B8",x"7E",x"DC",x"DA",x"5C",x"B7",x"7B",x"7D",x"D8",x"BF",x"AE",
x"AA",x"AB",x"DD",x"DE",x"DF",x"7F",x"B5",x"D6",x"7C",x"D5",x"5D",x"DB",x"B6",x"D9",x"5B",x"D7",
x"0C",x"07",x"06",x"04",x"05",x"08",x"0A",x"0B",x"09",x"0F",x"E2",x"2A",x"3F",x"CD",x"C8",x"CC",
x"CB",x"5E",x"AC",x"2D",x"2B",x"3D",x"2E",x"2C",x"3B",x"22",x"C7",x"3C",x"C3",x"3E",x"C5",x"2F",
x"C9",x"60",x"C6",x"3A",x"D0",x"CE",x"A8",x"CA",x"D3",x"D4",x"D1",x"D2",x"A9",x"CF",x"2E",x"2F",
x"11",x"FF",x"FF",x"01",x"FE",x"FE",x"ED",x"78",x"2F",x"E6",x"1F",x"28",x"0E",x"67",x"7D",x"14",
x"C0",x"D6",x"08",x"CB",x"3C",x"30",x"FA",x"53",x"5F",x"20",x"F4",x"2D",x"CB",x"00",x"38",x"E6",
x"7A",x"3C",x"C8",x"FE",x"28",x"C8",x"FE",x"19",x"C8",x"7B",x"5A",x"57",x"FE",x"18",x"C9",x"CD",
x"8E",x"02",x"C0",x"21",x"00",x"5C",x"CB",x"7E",x"20",x"07",x"23",x"35",x"2B",x"20",x"02",x"36",
x"FF",x"7D",x"21",x"04",x"5C",x"BD",x"20",x"EE",x"CD",x"1E",x"03",x"D0",x"21",x"00",x"5C",x"BE",
x"28",x"2E",x"EB",x"21",x"04",x"5C",x"BE",x"28",x"27",x"CB",x"7E",x"20",x"04",x"EB",x"CB",x"7E",
x"C8",x"5F",x"77",x"23",x"36",x"05",x"23",x"3A",x"09",x"5C",x"77",x"23",x"FD",x"4E",x"07",x"FD",
x"56",x"01",x"E5",x"CD",x"33",x"03",x"E1",x"77",x"32",x"08",x"5C",x"FD",x"CB",x"01",x"EE",x"C9",
x"23",x"36",x"05",x"23",x"35",x"C0",x"3A",x"0A",x"5C",x"77",x"23",x"7E",x"18",x"EA",x"42",x"16",
x"00",x"7B",x"FE",x"27",x"D0",x"FE",x"18",x"20",x"03",x"CB",x"78",x"C0",x"21",x"05",x"02",x"19",
x"7E",x"37",x"C9",x"7B",x"FE",x"3A",x"38",x"2F",x"0D",x"FA",x"4F",x"03",x"28",x"03",x"C6",x"4F",
x"C9",x"21",x"EB",x"01",x"04",x"28",x"03",x"21",x"05",x"02",x"16",x"00",x"19",x"7E",x"C9",x"21",
x"29",x"02",x"CB",x"40",x"28",x"F4",x"CB",x"5A",x"28",x"0A",x"FD",x"CB",x"30",x"5E",x"C0",x"04",
x"C0",x"C6",x"20",x"C9",x"C6",x"A5",x"C9",x"FE",x"30",x"D8",x"0D",x"FA",x"9D",x"03",x"20",x"19",
x"21",x"54",x"02",x"CB",x"68",x"28",x"D3",x"FE",x"38",x"30",x"07",x"D6",x"20",x"04",x"C8",x"C6",
x"08",x"C9",x"D6",x"36",x"04",x"C8",x"C6",x"FE",x"C9",x"21",x"30",x"02",x"FE",x"39",x"28",x"BA",
x"FE",x"30",x"28",x"B6",x"E6",x"07",x"C6",x"80",x"04",x"C8",x"EE",x"0F",x"C9",x"04",x"C8",x"CB",
x"68",x"21",x"30",x"02",x"20",x"A4",x"D6",x"10",x"FE",x"22",x"28",x"06",x"FE",x"20",x"C0",x"3E",
x"5F",x"C9",x"3E",x"40",x"C9",x"F3",x"7D",x"CB",x"3D",x"CB",x"3D",x"2F",x"E6",x"03",x"4F",x"06",
x"00",x"DD",x"21",x"D1",x"03",x"DD",x"09",x"3A",x"48",x"5C",x"E6",x"38",x"0F",x"0F",x"0F",x"F6",
x"08",x"00",x"00",x"00",x"04",x"0C",x"0D",x"20",x"FD",x"0E",x"3F",x"05",x"C2",x"D6",x"03",x"EE",
x"10",x"D3",x"FE",x"44",x"4F",x"CB",x"67",x"20",x"09",x"7A",x"B3",x"28",x"09",x"79",x"4D",x"1B",
x"DD",x"E9",x"4D",x"0C",x"DD",x"E9",x"FB",x"C9",x"EF",x"31",x"27",x"C0",x"03",x"34",x"EC",x"6C",
x"98",x"1F",x"F5",x"04",x"A1",x"0F",x"38",x"21",x"92",x"5C",x"7E",x"A7",x"20",x"5E",x"23",x"4E",
x"23",x"46",x"78",x"17",x"9F",x"B9",x"20",x"54",x"23",x"BE",x"20",x"50",x"78",x"C6",x"3C",x"F2",
x"25",x"04",x"E2",x"6C",x"04",x"06",x"FA",x"04",x"D6",x"0C",x"30",x"FB",x"C6",x"0C",x"C5",x"21",
x"6E",x"04",x"CD",x"06",x"34",x"CD",x"B4",x"33",x"EF",x"04",x"38",x"F1",x"86",x"77",x"EF",x"C0",
x"02",x"31",x"38",x"CD",x"94",x"1E",x"FE",x"0B",x"30",x"22",x"EF",x"E0",x"04",x"E0",x"34",x"80",
x"43",x"55",x"9F",x"80",x"01",x"05",x"34",x"35",x"71",x"03",x"38",x"CD",x"99",x"1E",x"C5",x"CD",
x"99",x"1E",x"E1",x"50",x"59",x"7A",x"B3",x"C8",x"1B",x"C3",x"B5",x"03",x"CF",x"0A",x"89",x"02",
x"D0",x"12",x"86",x"89",x"0A",x"97",x"60",x"75",x"89",x"12",x"D5",x"17",x"1F",x"89",x"1B",x"90",
x"41",x"02",x"89",x"24",x"D0",x"53",x"CA",x"89",x"2E",x"9D",x"36",x"B1",x"89",x"38",x"FF",x"49",
x"3E",x"89",x"43",x"FF",x"6A",x"73",x"89",x"4F",x"A7",x"00",x"54",x"89",x"5C",x"00",x"00",x"00",
x"89",x"69",x"14",x"F6",x"24",x"89",x"76",x"F1",x"10",x"05",x"CD",x"FB",x"24",x"3A",x"3B",x"5C",
x"87",x"FA",x"8A",x"1C",x"E1",x"D0",x"E5",x"CD",x"F1",x"2B",x"62",x"6B",x"0D",x"F8",x"09",x"CB",
x"FE",x"C9",x"21",x"3F",x"05",x"E5",x"21",x"80",x"1F",x"CB",x"7F",x"28",x"03",x"21",x"98",x"0C",
x"08",x"13",x"DD",x"2B",x"F3",x"3E",x"02",x"47",x"10",x"FE",x"D3",x"FE",x"EE",x"0F",x"06",x"A4",
x"2D",x"20",x"F5",x"05",x"25",x"F2",x"D8",x"04",x"06",x"2F",x"10",x"FE",x"D3",x"FE",x"3E",x"0D",
x"06",x"37",x"10",x"FE",x"D3",x"FE",x"01",x"0E",x"3B",x"08",x"6F",x"C3",x"07",x"05",x"7A",x"B3",
x"28",x"0C",x"DD",x"6E",x"00",x"7C",x"AD",x"67",x"3E",x"01",x"37",x"C3",x"25",x"05",x"6C",x"18",
x"F4",x"79",x"CB",x"78",x"10",x"FE",x"30",x"04",x"06",x"42",x"10",x"FE",x"D3",x"FE",x"06",x"3E",
x"20",x"EF",x"05",x"AF",x"3C",x"CB",x"15",x"C2",x"14",x"05",x"1B",x"DD",x"23",x"06",x"31",x"3E",
x"7F",x"DB",x"FE",x"1F",x"D0",x"7A",x"3C",x"C2",x"FE",x"04",x"06",x"3B",x"10",x"FE",x"C9",x"F5",
x"3A",x"48",x"5C",x"E6",x"38",x"0F",x"0F",x"0F",x"D3",x"FE",x"3E",x"7F",x"DB",x"FE",x"1F",x"FB",
x"38",x"02",x"CF",x"0C",x"F1",x"C9",x"F3",x"31",x"BF",x"04",x"DB",x"FB",x"ED",x"47",x"CD",x"DD",
x"05",x"E5",x"CD",x"DD",x"05",x"EB",x"CD",x"DD",x"05",x"44",x"4D",x"CD",x"DD",x"05",x"E5",x"F1",
x"08",x"E1",x"D9",x"CD",x"DD",x"05",x"22",x"B0",x"04",x"CD",x"DD",x"05",x"EB",x"CD",x"DD",x"05",
x"44",x"4D",x"CD",x"DD",x"05",x"E5",x"FD",x"E1",x"CD",x"DD",x"05",x"E5",x"DD",x"E1",x"DB",x"FB",
x"E6",x"02",x"0F",x"32",x"B2",x"04",x"DB",x"FB",x"ED",x"4F",x"CD",x"DD",x"05",x"E5",x"CD",x"DD",
x"05",x"22",x"B4",x"04",x"DB",x"FB",x"A7",x"28",x"07",x"3D",x"28",x"08",x"ED",x"5E",x"18",x"06",
x"ED",x"46",x"18",x"02",x"ED",x"56",x"DB",x"FB",x"E6",x"07",x"D3",x"FE",x"21",x"00",x"40",x"DB",
x"FB",x"77",x"23",x"7C",x"B5",x"20",x"F8",x"2A",x"B0",x"04",x"3A",x"B2",x"04",x"0F",x"38",x"06",
x"F1",x"ED",x"7B",x"B4",x"04",x"C9",x"F1",x"ED",x"7B",x"B4",x"04",x"FB",x"C9",x"DB",x"FB",x"6F",
x"DB",x"FB",x"67",x"C9",x"E7",x"05",x"D0",x"3E",x"16",x"3D",x"20",x"FD",x"A7",x"04",x"C8",x"3E",
x"7F",x"DB",x"FE",x"1F",x"D0",x"A9",x"E6",x"20",x"28",x"F3",x"79",x"2F",x"4F",x"E6",x"07",x"F6",
x"08",x"D3",x"FE",x"37",x"C9",x"F1",x"3A",x"74",x"5C",x"D6",x"E0",x"32",x"74",x"5C",x"CD",x"8C",
x"1C",x"CD",x"30",x"25",x"28",x"3C",x"01",x"11",x"00",x"3A",x"74",x"5C",x"A7",x"28",x"02",x"0E",
x"22",x"F7",x"D5",x"DD",x"E1",x"06",x"0B",x"3E",x"20",x"12",x"13",x"10",x"FC",x"DD",x"36",x"01",
x"FF",x"CD",x"F1",x"2B",x"21",x"F6",x"FF",x"0B",x"09",x"03",x"30",x"0F",x"3A",x"74",x"5C",x"A7",
x"20",x"02",x"CF",x"0E",x"78",x"B1",x"28",x"0A",x"01",x"0A",x"00",x"DD",x"E5",x"E1",x"23",x"EB",
x"ED",x"B0",x"DF",x"FE",x"E4",x"20",x"49",x"3A",x"74",x"5C",x"FE",x"03",x"CA",x"8A",x"1C",x"E7",
x"CD",x"B2",x"28",x"CB",x"F9",x"30",x"0B",x"21",x"00",x"00",x"3A",x"74",x"5C",x"3D",x"28",x"15",
x"CF",x"01",x"C2",x"8A",x"1C",x"CD",x"30",x"25",x"28",x"18",x"23",x"7E",x"DD",x"77",x"0B",x"23",
x"7E",x"DD",x"77",x"0C",x"23",x"DD",x"71",x"0E",x"3E",x"01",x"CB",x"71",x"28",x"01",x"3C",x"DD",
x"77",x"00",x"EB",x"E7",x"FE",x"29",x"20",x"DA",x"E7",x"CD",x"EE",x"1B",x"EB",x"C3",x"5A",x"07",
x"FE",x"AA",x"20",x"1F",x"3A",x"74",x"5C",x"FE",x"03",x"CA",x"8A",x"1C",x"E7",x"CD",x"EE",x"1B",
x"DD",x"36",x"0B",x"00",x"DD",x"36",x"0C",x"1B",x"21",x"00",x"40",x"DD",x"75",x"0D",x"DD",x"74",
x"0E",x"18",x"4D",x"FE",x"AF",x"20",x"4F",x"3A",x"74",x"5C",x"FE",x"03",x"CA",x"8A",x"1C",x"E7",
x"CD",x"48",x"20",x"20",x"0C",x"3A",x"74",x"5C",x"A7",x"CA",x"8A",x"1C",x"CD",x"E6",x"1C",x"18",
x"0F",x"CD",x"82",x"1C",x"DF",x"FE",x"2C",x"28",x"0C",x"3A",x"74",x"5C",x"A7",x"CA",x"8A",x"1C",
x"CD",x"E6",x"1C",x"18",x"04",x"E7",x"CD",x"82",x"1C",x"CD",x"EE",x"1B",x"CD",x"99",x"1E",x"DD",
x"71",x"0B",x"DD",x"70",x"0C",x"CD",x"99",x"1E",x"DD",x"71",x"0D",x"DD",x"70",x"0E",x"60",x"69",
x"DD",x"36",x"00",x"03",x"18",x"44",x"FE",x"CA",x"28",x"09",x"CD",x"EE",x"1B",x"DD",x"36",x"0E",
x"80",x"18",x"17",x"3A",x"74",x"5C",x"A7",x"C2",x"8A",x"1C",x"E7",x"CD",x"82",x"1C",x"CD",x"EE",
x"1B",x"CD",x"99",x"1E",x"DD",x"71",x"0D",x"DD",x"70",x"0E",x"DD",x"36",x"00",x"00",x"2A",x"59",
x"5C",x"ED",x"5B",x"53",x"5C",x"37",x"ED",x"52",x"DD",x"75",x"0B",x"DD",x"74",x"0C",x"2A",x"4B",
x"5C",x"ED",x"52",x"DD",x"75",x"0F",x"DD",x"74",x"10",x"EB",x"3A",x"74",x"5C",x"A7",x"CA",x"70",
x"09",x"E5",x"01",x"11",x"00",x"DD",x"09",x"DD",x"E5",x"11",x"11",x"00",x"AF",x"37",x"CD",x"56",
x"05",x"DD",x"E1",x"30",x"F2",x"3E",x"FE",x"CD",x"01",x"16",x"FD",x"36",x"52",x"03",x"0E",x"80",
x"DD",x"7E",x"00",x"DD",x"BE",x"EF",x"20",x"02",x"0E",x"F6",x"FE",x"04",x"30",x"D9",x"11",x"C0",
x"09",x"C5",x"CD",x"0A",x"0C",x"C1",x"DD",x"E5",x"D1",x"21",x"F0",x"FF",x"19",x"06",x"0A",x"7E",
x"3C",x"20",x"03",x"79",x"80",x"4F",x"13",x"1A",x"BE",x"23",x"20",x"01",x"0C",x"D7",x"10",x"F6",
x"CB",x"79",x"20",x"B3",x"3E",x"0D",x"D7",x"E1",x"DD",x"7E",x"00",x"FE",x"03",x"28",x"0C",x"3A",
x"74",x"5C",x"3D",x"CA",x"08",x"08",x"FE",x"02",x"CA",x"B6",x"08",x"E5",x"DD",x"6E",x"FA",x"DD",
x"66",x"FB",x"DD",x"5E",x"0B",x"DD",x"56",x"0C",x"7C",x"B5",x"28",x"0D",x"ED",x"52",x"38",x"26",
x"28",x"07",x"DD",x"7E",x"00",x"FE",x"03",x"20",x"1D",x"E1",x"7C",x"B5",x"20",x"06",x"DD",x"6E",
x"0D",x"DD",x"66",x"0E",x"E5",x"DD",x"E1",x"3A",x"74",x"5C",x"FE",x"02",x"37",x"20",x"01",x"A7",
x"3E",x"FF",x"CD",x"56",x"05",x"D8",x"CF",x"1A",x"DD",x"5E",x"0B",x"DD",x"56",x"0C",x"E5",x"7C",
x"B5",x"20",x"06",x"13",x"13",x"13",x"EB",x"18",x"0C",x"DD",x"6E",x"FA",x"DD",x"66",x"FB",x"EB",
x"37",x"ED",x"52",x"38",x"09",x"11",x"05",x"00",x"19",x"44",x"4D",x"CD",x"05",x"1F",x"E1",x"DD",
x"7E",x"00",x"A7",x"28",x"3E",x"7C",x"B5",x"28",x"13",x"2B",x"46",x"2B",x"4E",x"2B",x"03",x"03",
x"03",x"DD",x"22",x"5F",x"5C",x"CD",x"E8",x"19",x"DD",x"2A",x"5F",x"5C",x"2A",x"59",x"5C",x"2B",
x"DD",x"4E",x"0B",x"DD",x"46",x"0C",x"C5",x"03",x"03",x"03",x"DD",x"7E",x"FD",x"F5",x"CD",x"55",
x"16",x"23",x"F1",x"77",x"D1",x"23",x"73",x"23",x"72",x"23",x"E5",x"DD",x"E1",x"37",x"3E",x"FF",
x"C3",x"02",x"08",x"EB",x"2A",x"59",x"5C",x"2B",x"DD",x"22",x"5F",x"5C",x"DD",x"4E",x"0B",x"DD",
x"46",x"0C",x"C5",x"CD",x"E5",x"19",x"C1",x"E5",x"C5",x"CD",x"55",x"16",x"DD",x"2A",x"5F",x"5C",
x"23",x"DD",x"4E",x"0F",x"DD",x"46",x"10",x"09",x"22",x"4B",x"5C",x"DD",x"66",x"0E",x"7C",x"E6",
x"C0",x"20",x"0A",x"DD",x"6E",x"0D",x"22",x"42",x"5C",x"FD",x"36",x"0A",x"00",x"D1",x"DD",x"E1",
x"37",x"3E",x"FF",x"C3",x"02",x"08",x"DD",x"4E",x"0B",x"DD",x"46",x"0C",x"C5",x"03",x"F7",x"36",
x"80",x"EB",x"D1",x"E5",x"E5",x"DD",x"E1",x"37",x"3E",x"FF",x"CD",x"02",x"08",x"E1",x"ED",x"5B",
x"53",x"5C",x"7E",x"E6",x"C0",x"20",x"19",x"1A",x"13",x"BE",x"23",x"20",x"02",x"1A",x"BE",x"1B",
x"2B",x"30",x"08",x"E5",x"EB",x"CD",x"B8",x"19",x"E1",x"18",x"EC",x"CD",x"2C",x"09",x"18",x"E2",
x"7E",x"4F",x"FE",x"80",x"C8",x"E5",x"2A",x"4B",x"5C",x"7E",x"FE",x"80",x"28",x"25",x"B9",x"28",
x"08",x"C5",x"CD",x"B8",x"19",x"C1",x"EB",x"18",x"F0",x"E6",x"E0",x"FE",x"A0",x"20",x"12",x"D1",
x"D5",x"E5",x"23",x"13",x"1A",x"BE",x"20",x"06",x"17",x"30",x"F7",x"E1",x"18",x"03",x"E1",x"18",
x"E0",x"3E",x"FF",x"D1",x"EB",x"3C",x"37",x"CD",x"2C",x"09",x"18",x"C4",x"20",x"10",x"08",x"22",
x"5F",x"5C",x"EB",x"CD",x"B8",x"19",x"CD",x"E8",x"19",x"EB",x"2A",x"5F",x"5C",x"08",x"08",x"D5",
x"CD",x"B8",x"19",x"22",x"5F",x"5C",x"2A",x"53",x"5C",x"E3",x"C5",x"08",x"38",x"07",x"2B",x"CD",
x"55",x"16",x"23",x"18",x"03",x"CD",x"55",x"16",x"23",x"C1",x"D1",x"ED",x"53",x"53",x"5C",x"ED",
x"5B",x"5F",x"5C",x"C5",x"D5",x"EB",x"ED",x"B0",x"E1",x"C1",x"D5",x"CD",x"E8",x"19",x"D1",x"C9",
x"E5",x"3E",x"FD",x"CD",x"01",x"16",x"AF",x"11",x"A1",x"09",x"CD",x"0A",x"0C",x"FD",x"CB",x"02",
x"EE",x"CD",x"D4",x"15",x"DD",x"E5",x"11",x"11",x"00",x"AF",x"CD",x"C2",x"04",x"DD",x"E1",x"06",
x"32",x"76",x"10",x"FD",x"DD",x"5E",x"0B",x"DD",x"56",x"0C",x"3E",x"FF",x"DD",x"E1",x"C3",x"C2",
x"04",x"80",x"53",x"74",x"61",x"72",x"74",x"20",x"74",x"61",x"70",x"65",x"2C",x"20",x"74",x"68",
x"65",x"6E",x"20",x"70",x"72",x"65",x"73",x"73",x"20",x"61",x"6E",x"79",x"20",x"6B",x"65",x"79",
x"AE",x"0D",x"50",x"72",x"6F",x"67",x"72",x"61",x"6D",x"3A",x"A0",x"0D",x"4E",x"75",x"6D",x"62",
x"65",x"72",x"20",x"61",x"72",x"72",x"61",x"79",x"3A",x"A0",x"0D",x"43",x"68",x"61",x"72",x"61",
x"63",x"74",x"65",x"72",x"20",x"61",x"72",x"72",x"61",x"79",x"3A",x"A0",x"0D",x"42",x"79",x"74",
x"65",x"73",x"3A",x"A0",x"CD",x"03",x"0B",x"FE",x"20",x"D2",x"D9",x"0A",x"FE",x"06",x"38",x"69",
x"FE",x"18",x"30",x"65",x"21",x"0B",x"0A",x"5F",x"16",x"00",x"19",x"5E",x"19",x"E5",x"C3",x"03",
x"0B",x"4E",x"57",x"10",x"29",x"54",x"53",x"52",x"37",x"50",x"4F",x"5F",x"5E",x"5D",x"5C",x"5B",
x"5A",x"54",x"53",x"0C",x"3E",x"22",x"B9",x"20",x"11",x"FD",x"CB",x"01",x"4E",x"20",x"09",x"04",
x"0E",x"02",x"3E",x"18",x"B8",x"20",x"03",x"05",x"0E",x"21",x"C3",x"D9",x"0D",x"3A",x"91",x"5C",
x"F5",x"FD",x"36",x"57",x"01",x"3E",x"20",x"CD",x"65",x"0B",x"F1",x"32",x"91",x"5C",x"C9",x"FD",
x"CB",x"01",x"4E",x"C2",x"CD",x"0E",x"0E",x"21",x"CD",x"55",x"0C",x"05",x"C3",x"D9",x"0D",x"CD",
x"03",x"0B",x"79",x"3D",x"3D",x"E6",x"10",x"18",x"5A",x"3E",x"3F",x"18",x"6C",x"11",x"87",x"0A",
x"32",x"0F",x"5C",x"18",x"0B",x"11",x"6D",x"0A",x"18",x"03",x"11",x"87",x"0A",x"32",x"0E",x"5C",
x"2A",x"51",x"5C",x"73",x"23",x"72",x"C9",x"11",x"F4",x"09",x"CD",x"80",x"0A",x"2A",x"0E",x"5C",
x"57",x"7D",x"FE",x"16",x"DA",x"11",x"22",x"20",x"29",x"44",x"4A",x"3E",x"1F",x"91",x"38",x"0C",
x"C6",x"02",x"4F",x"FD",x"CB",x"01",x"4E",x"20",x"16",x"3E",x"16",x"90",x"DA",x"9F",x"1E",x"3C",
x"47",x"04",x"FD",x"CB",x"02",x"46",x"C2",x"55",x"0C",x"FD",x"BE",x"31",x"DA",x"86",x"0C",x"C3",
x"D9",x"0D",x"7C",x"CD",x"03",x"0B",x"81",x"3D",x"E6",x"1F",x"C8",x"57",x"FD",x"CB",x"01",x"C6",
x"3E",x"20",x"CD",x"3B",x"0C",x"15",x"20",x"F8",x"C9",x"CD",x"24",x"0B",x"FD",x"CB",x"01",x"4E",
x"20",x"1A",x"FD",x"CB",x"02",x"46",x"20",x"08",x"ED",x"43",x"88",x"5C",x"22",x"84",x"5C",x"C9",
x"ED",x"43",x"8A",x"5C",x"ED",x"43",x"82",x"5C",x"22",x"86",x"5C",x"C9",x"FD",x"71",x"45",x"22",
x"80",x"5C",x"C9",x"FD",x"CB",x"01",x"4E",x"20",x"14",x"ED",x"4B",x"88",x"5C",x"2A",x"84",x"5C",
x"FD",x"CB",x"02",x"46",x"C8",x"ED",x"4B",x"8A",x"5C",x"2A",x"86",x"5C",x"C9",x"FD",x"4E",x"45",
x"2A",x"80",x"5C",x"C9",x"FE",x"80",x"38",x"3D",x"FE",x"90",x"30",x"26",x"47",x"CD",x"38",x"0B",
x"CD",x"03",x"0B",x"11",x"92",x"5C",x"18",x"47",x"21",x"92",x"5C",x"CD",x"3E",x"0B",x"CB",x"18",
x"9F",x"E6",x"0F",x"4F",x"CB",x"18",x"9F",x"E6",x"F0",x"B1",x"0E",x"04",x"77",x"23",x"0D",x"20",
x"FB",x"C9",x"D6",x"A5",x"30",x"09",x"C6",x"15",x"C5",x"ED",x"4B",x"7B",x"5C",x"18",x"0B",x"CD",
x"10",x"0C",x"C3",x"03",x"0B",x"C5",x"ED",x"4B",x"36",x"5C",x"EB",x"21",x"3B",x"5C",x"CB",x"86",
x"FE",x"20",x"20",x"02",x"CB",x"C6",x"26",x"00",x"6F",x"29",x"29",x"29",x"09",x"C1",x"EB",x"79",
x"3D",x"3E",x"21",x"20",x"0E",x"05",x"4F",x"FD",x"CB",x"01",x"4E",x"28",x"06",x"D5",x"CD",x"CD",
x"0E",x"D1",x"79",x"B9",x"D5",x"CC",x"55",x"0C",x"D1",x"C5",x"E5",x"3A",x"91",x"5C",x"06",x"FF",
x"1F",x"38",x"01",x"04",x"1F",x"1F",x"9F",x"4F",x"3E",x"08",x"A7",x"FD",x"CB",x"01",x"4E",x"28",
x"05",x"FD",x"CB",x"30",x"CE",x"37",x"EB",x"08",x"1A",x"A0",x"AE",x"A9",x"12",x"08",x"38",x"13",
x"14",x"23",x"3D",x"20",x"F2",x"EB",x"25",x"FD",x"CB",x"01",x"4E",x"CC",x"DB",x"0B",x"E1",x"C1",
x"0D",x"23",x"C9",x"08",x"3E",x"20",x"83",x"5F",x"08",x"18",x"E6",x"7C",x"0F",x"0F",x"0F",x"E6",
x"03",x"F6",x"58",x"67",x"ED",x"5B",x"8F",x"5C",x"7E",x"AB",x"A2",x"AB",x"FD",x"CB",x"57",x"76",
x"28",x"08",x"E6",x"C7",x"CB",x"57",x"20",x"02",x"EE",x"38",x"FD",x"CB",x"57",x"66",x"28",x"08",
x"E6",x"F8",x"CB",x"6F",x"20",x"02",x"EE",x"07",x"77",x"C9",x"E5",x"26",x"00",x"E3",x"18",x"04",
x"11",x"95",x"00",x"F5",x"CD",x"41",x"0C",x"38",x"09",x"3E",x"20",x"FD",x"CB",x"01",x"46",x"CC",
x"3B",x"0C",x"1A",x"E6",x"7F",x"CD",x"3B",x"0C",x"1A",x"13",x"87",x"30",x"F5",x"D1",x"FE",x"48",
x"28",x"03",x"FE",x"82",x"D8",x"7A",x"FE",x"03",x"D8",x"3E",x"20",x"D5",x"D9",x"D7",x"D9",x"D1",
x"C9",x"F5",x"EB",x"3C",x"CB",x"7E",x"23",x"28",x"FB",x"3D",x"20",x"F8",x"EB",x"F1",x"FE",x"20",
x"D8",x"1A",x"D6",x"41",x"C9",x"FD",x"CB",x"01",x"4E",x"C0",x"11",x"D9",x"0D",x"D5",x"78",x"FD",
x"CB",x"02",x"46",x"C2",x"02",x"0D",x"FD",x"BE",x"31",x"38",x"1B",x"C0",x"FD",x"CB",x"02",x"66",
x"28",x"16",x"FD",x"5E",x"2D",x"1D",x"28",x"5A",x"3E",x"00",x"CD",x"01",x"16",x"ED",x"7B",x"3F",
x"5C",x"FD",x"CB",x"02",x"A6",x"C9",x"CF",x"04",x"FD",x"35",x"52",x"20",x"45",x"3E",x"18",x"90",
x"32",x"8C",x"5C",x"2A",x"8F",x"5C",x"E5",x"3A",x"91",x"5C",x"F5",x"3E",x"FD",x"CD",x"01",x"16",
x"AF",x"11",x"F8",x"0C",x"CD",x"0A",x"0C",x"FD",x"CB",x"02",x"EE",x"21",x"3B",x"5C",x"CB",x"DE",
x"CB",x"AE",x"D9",x"CD",x"D4",x"15",x"D9",x"FE",x"20",x"CA",x"77",x"38",x"FE",x"E2",x"CA",x"77",
x"38",x"C3",x"70",x"38",x"00",x"3E",x"FE",x"CD",x"01",x"16",x"F1",x"32",x"91",x"5C",x"E1",x"22",
x"8F",x"5C",x"CD",x"FE",x"0D",x"FD",x"46",x"31",x"04",x"0E",x"21",x"C5",x"CD",x"9B",x"0E",x"7C",
x"0F",x"0F",x"0F",x"E6",x"03",x"F6",x"58",x"67",x"11",x"E0",x"5A",x"1A",x"4E",x"06",x"20",x"EB",
x"12",x"71",x"13",x"23",x"10",x"FA",x"C1",x"C9",x"80",x"73",x"63",x"72",x"6F",x"6C",x"6C",x"BF",
x"CF",x"0C",x"FE",x"02",x"38",x"80",x"FD",x"86",x"31",x"D6",x"19",x"D0",x"ED",x"44",x"C5",x"47",
x"2A",x"8F",x"5C",x"E5",x"2A",x"91",x"5C",x"E5",x"CD",x"4D",x"0D",x"78",x"F5",x"21",x"6B",x"5C",
x"46",x"78",x"3C",x"77",x"21",x"89",x"5C",x"BE",x"38",x"03",x"34",x"06",x"18",x"CD",x"00",x"0E",
x"F1",x"3D",x"20",x"E8",x"E1",x"FD",x"75",x"57",x"E1",x"22",x"8F",x"5C",x"ED",x"4B",x"88",x"5C",
x"FD",x"CB",x"02",x"86",x"CD",x"D9",x"0D",x"FD",x"CB",x"02",x"C6",x"C1",x"C9",x"AF",x"2A",x"8D",
x"5C",x"FD",x"CB",x"02",x"46",x"28",x"04",x"67",x"FD",x"6E",x"0E",x"22",x"8F",x"5C",x"21",x"91",
x"5C",x"20",x"02",x"7E",x"0F",x"AE",x"E6",x"55",x"AE",x"77",x"C9",x"CD",x"AF",x"0D",x"21",x"3C",
x"5C",x"CB",x"AE",x"CB",x"C6",x"CD",x"4D",x"0D",x"FD",x"46",x"31",x"CD",x"44",x"0E",x"21",x"C0",
x"5A",x"3A",x"8D",x"5C",x"05",x"18",x"07",x"0E",x"20",x"2B",x"77",x"0D",x"20",x"FB",x"10",x"F7",
x"FD",x"36",x"31",x"02",x"3E",x"FD",x"CD",x"01",x"16",x"2A",x"51",x"5C",x"11",x"F4",x"09",x"A7",
x"73",x"23",x"72",x"23",x"11",x"A8",x"10",x"3F",x"38",x"F6",x"01",x"21",x"17",x"18",x"2A",x"21",
x"00",x"00",x"22",x"7D",x"5C",x"FD",x"CB",x"30",x"86",x"CD",x"94",x"0D",x"3E",x"FE",x"CD",x"01",
x"16",x"CD",x"4D",x"0D",x"06",x"18",x"CD",x"44",x"0E",x"2A",x"51",x"5C",x"11",x"F4",x"09",x"73",
x"23",x"72",x"FD",x"36",x"52",x"01",x"01",x"21",x"18",x"21",x"00",x"5B",x"FD",x"CB",x"01",x"4E",
x"20",x"12",x"78",x"FD",x"CB",x"02",x"46",x"28",x"05",x"FD",x"86",x"31",x"D6",x"18",x"C5",x"47",
x"CD",x"9B",x"0E",x"C1",x"3E",x"21",x"91",x"5F",x"16",x"00",x"19",x"C3",x"DC",x"0A",x"06",x"17",
x"CD",x"9B",x"0E",x"0E",x"08",x"C5",x"E5",x"78",x"E6",x"07",x"78",x"20",x"0C",x"EB",x"21",x"E0",
x"F8",x"19",x"EB",x"01",x"20",x"00",x"3D",x"ED",x"B0",x"EB",x"21",x"E0",x"FF",x"19",x"EB",x"47",
x"E6",x"07",x"0F",x"0F",x"0F",x"4F",x"78",x"06",x"00",x"ED",x"B0",x"06",x"07",x"09",x"E6",x"F8",
x"20",x"DB",x"E1",x"24",x"C1",x"0D",x"20",x"CD",x"CD",x"88",x"0E",x"21",x"E0",x"FF",x"19",x"EB",
x"ED",x"B0",x"06",x"01",x"C5",x"CD",x"9B",x"0E",x"0E",x"08",x"C5",x"E5",x"78",x"E6",x"07",x"0F",
x"0F",x"0F",x"4F",x"78",x"06",x"00",x"0D",x"54",x"5D",x"36",x"00",x"13",x"ED",x"B0",x"11",x"01",
x"07",x"19",x"3D",x"E6",x"F8",x"47",x"20",x"E5",x"E1",x"24",x"C1",x"0D",x"20",x"DC",x"CD",x"88",
x"0E",x"62",x"6B",x"13",x"3A",x"8D",x"5C",x"FD",x"CB",x"02",x"46",x"28",x"03",x"3A",x"48",x"5C",
x"77",x"0B",x"ED",x"B0",x"C1",x"0E",x"21",x"C9",x"7C",x"0F",x"0F",x"0F",x"3D",x"F6",x"50",x"67",
x"EB",x"61",x"68",x"29",x"29",x"29",x"29",x"29",x"44",x"4D",x"C9",x"3E",x"18",x"90",x"57",x"0F",
x"0F",x"0F",x"E6",x"E0",x"6F",x"7A",x"E6",x"18",x"F6",x"40",x"67",x"C9",x"CD",x"30",x"25",x"CA",
x"B2",x"1B",x"C3",x"91",x"38",x"3E",x"FF",x"D3",x"F7",x"DB",x"EF",x"0F",x"38",x"FB",x"DB",x"F7",
x"C9",x"20",x"6F",x"3F",x"9F",x"E6",x"F8",x"84",x"67",x"10",x"E7",x"18",x"0D",x"F3",x"21",x"00",
x"5B",x"06",x"08",x"C5",x"CD",x"F4",x"0E",x"C1",x"10",x"F9",x"3E",x"04",x"D3",x"FB",x"FB",x"21",
x"00",x"5B",x"FD",x"75",x"46",x"AF",x"47",x"77",x"23",x"10",x"FC",x"FD",x"CB",x"30",x"8E",x"0E",
x"21",x"C3",x"D9",x"0D",x"78",x"FE",x"03",x"9F",x"E6",x"02",x"D3",x"FB",x"57",x"CD",x"54",x"1F",
x"38",x"0A",x"3E",x"04",x"D3",x"FB",x"FB",x"CD",x"DF",x"0E",x"CF",x"0C",x"DB",x"FB",x"87",x"F8",
x"30",x"EB",x"0E",x"20",x"5E",x"23",x"06",x"08",x"CB",x"12",x"CB",x"13",x"CB",x"1A",x"DB",x"FB",
x"1F",x"30",x"FB",x"7A",x"D3",x"FB",x"10",x"F0",x"0D",x"20",x"E9",x"C9",x"2A",x"3D",x"5C",x"E5",
x"21",x"7F",x"10",x"E5",x"ED",x"73",x"3D",x"5C",x"CD",x"D4",x"15",x"F5",x"16",x"00",x"FD",x"5E",
x"FF",x"21",x"C8",x"00",x"CD",x"B5",x"03",x"F1",x"21",x"38",x"0F",x"E5",x"FE",x"18",x"30",x"31",
x"FE",x"07",x"38",x"2D",x"FE",x"10",x"38",x"3A",x"01",x"02",x"00",x"57",x"FE",x"16",x"38",x"0C",
x"03",x"FD",x"CB",x"37",x"7E",x"CA",x"1E",x"10",x"CD",x"D4",x"15",x"5F",x"CD",x"D4",x"15",x"D5",
x"2A",x"5B",x"5C",x"FD",x"CB",x"07",x"86",x"CD",x"55",x"16",x"C1",x"23",x"70",x"23",x"71",x"18",
x"0A",x"FD",x"CB",x"07",x"86",x"2A",x"5B",x"5C",x"CD",x"52",x"16",x"12",x"13",x"ED",x"53",x"5B",
x"5C",x"C9",x"5F",x"16",x"00",x"21",x"99",x"0F",x"19",x"5E",x"19",x"E5",x"2A",x"5B",x"5C",x"C9",
x"09",x"66",x"6A",x"50",x"B5",x"70",x"7E",x"CF",x"D4",x"2A",x"49",x"5C",x"FD",x"CB",x"37",x"6E",
x"C2",x"97",x"10",x"CD",x"6E",x"19",x"CD",x"95",x"16",x"7A",x"B3",x"CA",x"97",x"10",x"E5",x"23",
x"4E",x"23",x"46",x"21",x"0A",x"00",x"09",x"44",x"4D",x"CD",x"05",x"1F",x"CD",x"97",x"10",x"2A",
x"51",x"5C",x"E3",x"E5",x"3E",x"FF",x"CD",x"01",x"16",x"E1",x"2B",x"FD",x"35",x"0F",x"CD",x"55",
x"18",x"FD",x"34",x"0F",x"2A",x"59",x"5C",x"23",x"23",x"23",x"23",x"22",x"5B",x"5C",x"E1",x"CD",
x"15",x"16",x"C9",x"FD",x"CB",x"37",x"6E",x"20",x"08",x"21",x"49",x"5C",x"CD",x"0F",x"19",x"18",
x"6D",x"FD",x"36",x"00",x"10",x"18",x"1D",x"CD",x"31",x"10",x"18",x"05",x"7E",x"FE",x"0D",x"C8",
x"23",x"22",x"5B",x"5C",x"C9",x"CD",x"31",x"10",x"01",x"01",x"00",x"C3",x"E8",x"19",x"CD",x"D4",
x"15",x"CD",x"D4",x"15",x"E1",x"E1",x"E1",x"22",x"3D",x"5C",x"FD",x"CB",x"00",x"7E",x"C0",x"F9",
x"C9",x"37",x"CD",x"95",x"11",x"ED",x"52",x"19",x"23",x"C1",x"D8",x"C5",x"44",x"4D",x"62",x"6B",
x"23",x"1A",x"E6",x"F0",x"FE",x"10",x"20",x"09",x"23",x"1A",x"D6",x"17",x"CE",x"00",x"20",x"01",
x"23",x"A7",x"ED",x"42",x"09",x"EB",x"38",x"E6",x"C9",x"FD",x"CB",x"37",x"6E",x"C0",x"2A",x"49",
x"5C",x"CD",x"6E",x"19",x"EB",x"CD",x"95",x"16",x"21",x"4A",x"5C",x"CD",x"1C",x"19",x"CD",x"95",
x"17",x"3E",x"00",x"C3",x"01",x"16",x"FD",x"CB",x"37",x"7E",x"28",x"A8",x"C3",x"81",x"0F",x"FD",
x"CB",x"30",x"66",x"28",x"A1",x"FD",x"36",x"00",x"FF",x"16",x"00",x"FD",x"5E",x"FE",x"21",x"90",
x"1A",x"CD",x"B5",x"03",x"C3",x"30",x"0F",x"E5",x"CD",x"90",x"11",x"2B",x"CD",x"E5",x"19",x"22",
x"5B",x"5C",x"FD",x"36",x"07",x"00",x"E1",x"C9",x"FD",x"CB",x"02",x"5E",x"C4",x"1D",x"11",x"A7",
x"FD",x"CB",x"01",x"6E",x"C8",x"3A",x"08",x"5C",x"FD",x"CB",x"01",x"AE",x"F5",x"FD",x"CB",x"02",
x"6E",x"C4",x"6E",x"0D",x"F1",x"FE",x"20",x"30",x"52",x"FE",x"10",x"30",x"2D",x"FE",x"06",x"30",
x"0A",x"47",x"E6",x"01",x"4F",x"78",x"1F",x"C6",x"12",x"18",x"2A",x"20",x"09",x"21",x"6A",x"5C",
x"3E",x"08",x"AE",x"77",x"18",x"0E",x"FE",x"0E",x"D8",x"D6",x"0D",x"21",x"41",x"5C",x"BE",x"77",
x"20",x"02",x"36",x"00",x"FD",x"CB",x"02",x"DE",x"BF",x"C9",x"47",x"E6",x"07",x"4F",x"3E",x"10",
x"CB",x"58",x"20",x"01",x"3C",x"FD",x"71",x"D3",x"11",x"0D",x"11",x"18",x"06",x"3A",x"0D",x"5C",
x"11",x"A8",x"10",x"2A",x"4F",x"5C",x"23",x"23",x"73",x"23",x"72",x"37",x"C9",x"CD",x"4D",x"0D",
x"FD",x"CB",x"02",x"9E",x"FD",x"CB",x"02",x"AE",x"2A",x"8A",x"5C",x"E5",x"2A",x"3D",x"5C",x"E5",
x"21",x"67",x"11",x"E5",x"ED",x"73",x"3D",x"5C",x"2A",x"82",x"5C",x"E5",x"37",x"CD",x"95",x"11",
x"EB",x"CD",x"7D",x"18",x"EB",x"CD",x"E1",x"18",x"2A",x"8A",x"5C",x"E3",x"EB",x"CD",x"4D",x"0D",
x"3A",x"8B",x"5C",x"92",x"38",x"26",x"20",x"06",x"7B",x"FD",x"96",x"50",x"30",x"1E",x"3E",x"20",
x"D5",x"CD",x"F4",x"09",x"D1",x"18",x"E9",x"16",x"00",x"FD",x"5E",x"FE",x"21",x"90",x"1A",x"CD",
x"B5",x"03",x"FD",x"36",x"00",x"FF",x"ED",x"5B",x"8A",x"5C",x"18",x"02",x"D1",x"E1",x"E1",x"22",
x"3D",x"5C",x"C1",x"D5",x"CD",x"D9",x"0D",x"E1",x"22",x"82",x"5C",x"FD",x"36",x"26",x"00",x"C9",
x"2A",x"61",x"5C",x"2B",x"A7",x"ED",x"5B",x"59",x"5C",x"FD",x"CB",x"37",x"6E",x"C8",x"ED",x"5B",
x"61",x"5C",x"D8",x"2A",x"63",x"5C",x"C9",x"7E",x"FE",x"0E",x"01",x"06",x"00",x"CC",x"E8",x"19",
x"7E",x"23",x"FE",x"0D",x"20",x"F1",x"C9",x"F3",x"3E",x"FF",x"ED",x"5B",x"B2",x"5C",x"D9",x"ED",
x"4B",x"B4",x"5C",x"ED",x"5B",x"38",x"5C",x"2A",x"7B",x"5C",x"D9",x"47",x"3E",x"07",x"D3",x"FE",
x"3E",x"3F",x"ED",x"47",x"00",x"00",x"00",x"00",x"00",x"00",x"62",x"6B",x"36",x"02",x"2B",x"BC",
x"20",x"FA",x"A7",x"ED",x"52",x"19",x"23",x"30",x"06",x"35",x"28",x"03",x"35",x"28",x"F3",x"2B",
x"D9",x"ED",x"43",x"B4",x"5C",x"ED",x"53",x"38",x"5C",x"22",x"7B",x"5C",x"D9",x"04",x"28",x"19",
x"22",x"B4",x"5C",x"11",x"AF",x"3E",x"01",x"A8",x"00",x"EB",x"ED",x"B8",x"EB",x"23",x"22",x"7B",
x"5C",x"2B",x"01",x"40",x"00",x"ED",x"43",x"38",x"5C",x"22",x"B2",x"5C",x"21",x"00",x"3C",x"22",
x"36",x"5C",x"2A",x"B2",x"5C",x"36",x"3E",x"2B",x"F9",x"2B",x"2B",x"22",x"3D",x"5C",x"ED",x"56",
x"FD",x"21",x"3A",x"5C",x"FB",x"21",x"B6",x"5C",x"22",x"4F",x"5C",x"11",x"AF",x"15",x"01",x"15",
x"00",x"EB",x"ED",x"B0",x"EB",x"2B",x"22",x"57",x"5C",x"23",x"22",x"53",x"5C",x"22",x"4B",x"5C",
x"36",x"80",x"23",x"22",x"59",x"5C",x"36",x"0D",x"23",x"36",x"80",x"23",x"22",x"61",x"5C",x"22",
x"63",x"5C",x"22",x"65",x"5C",x"3E",x"38",x"32",x"8D",x"5C",x"32",x"8F",x"5C",x"32",x"48",x"5C",
x"21",x"23",x"05",x"22",x"09",x"5C",x"FD",x"35",x"C6",x"FD",x"35",x"CA",x"21",x"C6",x"15",x"11",
x"10",x"5C",x"01",x"0E",x"00",x"ED",x"B0",x"FD",x"CB",x"01",x"CE",x"CD",x"DF",x"0E",x"FD",x"36",
x"31",x"02",x"CD",x"6B",x"0D",x"AF",x"11",x"38",x"15",x"CD",x"0A",x"0C",x"FD",x"CB",x"02",x"EE",
x"18",x"07",x"FD",x"36",x"31",x"02",x"CD",x"95",x"17",x"CD",x"B0",x"16",x"3E",x"00",x"CD",x"01",
x"16",x"CD",x"2C",x"0F",x"CD",x"17",x"1B",x"FD",x"CB",x"00",x"7E",x"20",x"12",x"FD",x"CB",x"30",
x"66",x"28",x"40",x"2A",x"59",x"5C",x"CD",x"A7",x"11",x"FD",x"36",x"00",x"FF",x"18",x"DD",x"2A",
x"59",x"5C",x"22",x"5D",x"5C",x"CD",x"FB",x"19",x"78",x"B1",x"C2",x"5D",x"15",x"DF",x"FE",x"0D",
x"28",x"C0",x"FD",x"CB",x"30",x"46",x"C4",x"AF",x"0D",x"CD",x"6E",x"0D",x"3E",x"19",x"FD",x"96",
x"4F",x"32",x"8C",x"5C",x"FD",x"CB",x"01",x"FE",x"FD",x"36",x"00",x"FF",x"FD",x"36",x"0A",x"01",
x"CD",x"8A",x"1B",x"76",x"FD",x"CB",x"01",x"AE",x"FD",x"CB",x"30",x"4E",x"C4",x"CD",x"0E",x"3A",
x"3A",x"5C",x"3C",x"F5",x"21",x"00",x"00",x"FD",x"74",x"37",x"FD",x"74",x"26",x"22",x"0B",x"5C",
x"21",x"01",x"00",x"22",x"16",x"5C",x"CD",x"B0",x"16",x"FD",x"CB",x"37",x"AE",x"CD",x"6E",x"0D",
x"FD",x"CB",x"02",x"EE",x"F1",x"47",x"FE",x"0A",x"38",x"02",x"C6",x"07",x"CD",x"EF",x"15",x"3E",
x"20",x"D7",x"78",x"11",x"91",x"13",x"CD",x"0A",x"0C",x"AF",x"11",x"36",x"15",x"CD",x"0A",x"0C",
x"ED",x"4B",x"45",x"5C",x"CD",x"1B",x"1A",x"3E",x"3A",x"D7",x"FD",x"4E",x"0D",x"06",x"00",x"CD",
x"1B",x"1A",x"CD",x"97",x"10",x"3A",x"3A",x"5C",x"3C",x"28",x"1B",x"FE",x"09",x"28",x"04",x"FE",
x"15",x"20",x"03",x"FD",x"34",x"0D",x"01",x"03",x"00",x"11",x"70",x"5C",x"21",x"44",x"5C",x"CB",
x"7E",x"28",x"01",x"09",x"ED",x"B8",x"FD",x"36",x"0A",x"FF",x"FD",x"CB",x"01",x"9E",x"C3",x"AC",
x"12",x"80",x"4F",x"CB",x"4E",x"45",x"58",x"54",x"20",x"77",x"69",x"74",x"68",x"6F",x"75",x"74",
x"20",x"46",x"4F",x"D2",x"56",x"61",x"72",x"69",x"61",x"62",x"6C",x"65",x"20",x"6E",x"6F",x"74",
x"20",x"66",x"6F",x"75",x"6E",x"E4",x"53",x"75",x"62",x"73",x"63",x"72",x"69",x"70",x"74",x"20",
x"77",x"72",x"6F",x"6E",x"E7",x"4F",x"75",x"74",x"20",x"6F",x"66",x"20",x"6D",x"65",x"6D",x"6F",
x"72",x"F9",x"4F",x"75",x"74",x"20",x"6F",x"66",x"20",x"73",x"63",x"72",x"65",x"65",x"EE",x"4E",
x"75",x"6D",x"62",x"65",x"72",x"20",x"74",x"6F",x"6F",x"20",x"62",x"69",x"E7",x"52",x"45",x"54",
x"55",x"52",x"4E",x"20",x"77",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",x"47",x"4F",x"53",x"55",
x"C2",x"45",x"6E",x"64",x"20",x"6F",x"66",x"20",x"66",x"69",x"6C",x"E5",x"53",x"54",x"4F",x"50",
x"20",x"73",x"74",x"61",x"74",x"65",x"6D",x"65",x"6E",x"F4",x"49",x"6E",x"76",x"61",x"6C",x"69",
x"64",x"20",x"61",x"72",x"67",x"75",x"6D",x"65",x"6E",x"F4",x"49",x"6E",x"74",x"65",x"67",x"65",
x"72",x"20",x"6F",x"75",x"74",x"20",x"6F",x"66",x"20",x"72",x"61",x"6E",x"67",x"E5",x"4E",x"6F",
x"6E",x"73",x"65",x"6E",x"73",x"65",x"20",x"69",x"6E",x"20",x"42",x"41",x"53",x"49",x"C3",x"42",
x"52",x"45",x"41",x"4B",x"20",x"2D",x"20",x"43",x"4F",x"4E",x"54",x"20",x"72",x"65",x"70",x"65",
x"61",x"74",x"F3",x"4F",x"75",x"74",x"20",x"6F",x"66",x"20",x"44",x"41",x"54",x"C1",x"49",x"6E",
x"76",x"61",x"6C",x"69",x"64",x"20",x"66",x"69",x"6C",x"65",x"20",x"6E",x"61",x"6D",x"E5",x"4E",
x"6F",x"20",x"72",x"6F",x"6F",x"6D",x"20",x"66",x"6F",x"72",x"20",x"6C",x"69",x"6E",x"E5",x"53",
x"54",x"4F",x"50",x"20",x"69",x"6E",x"20",x"49",x"4E",x"50",x"55",x"D4",x"46",x"4F",x"52",x"20",
x"77",x"69",x"74",x"68",x"6F",x"75",x"74",x"20",x"4E",x"45",x"58",x"D4",x"49",x"6E",x"76",x"61",
x"6C",x"69",x"64",x"20",x"49",x"2F",x"4F",x"20",x"64",x"65",x"76",x"69",x"63",x"E5",x"49",x"6E",
x"76",x"61",x"6C",x"69",x"64",x"20",x"63",x"6F",x"6C",x"6F",x"75",x"F2",x"42",x"52",x"45",x"41",
x"4B",x"20",x"69",x"6E",x"74",x"6F",x"20",x"70",x"72",x"6F",x"67",x"72",x"61",x"ED",x"52",x"41",
x"4D",x"54",x"4F",x"50",x"20",x"6E",x"6F",x"20",x"67",x"6F",x"6F",x"E4",x"53",x"74",x"61",x"74",
x"65",x"6D",x"65",x"6E",x"74",x"20",x"6C",x"6F",x"73",x"F4",x"49",x"6E",x"76",x"61",x"6C",x"69",
x"64",x"20",x"73",x"74",x"72",x"65",x"61",x"ED",x"46",x"4E",x"20",x"77",x"69",x"74",x"68",x"6F",
x"75",x"74",x"20",x"44",x"45",x"C6",x"50",x"61",x"72",x"61",x"6D",x"65",x"74",x"65",x"72",x"20",
x"65",x"72",x"72",x"6F",x"F2",x"54",x"61",x"70",x"65",x"20",x"6C",x"6F",x"61",x"64",x"69",x"6E",
x"67",x"20",x"65",x"72",x"72",x"6F",x"F2",x"2C",x"A0",x"7F",x"20",x"31",x"39",x"38",x"32",x"20",
x"53",x"69",x"6E",x"63",x"6C",x"61",x"69",x"72",x"20",x"52",x"65",x"73",x"65",x"61",x"72",x"63",
x"68",x"20",x"4C",x"74",x"E4",x"3E",x"10",x"01",x"00",x"00",x"C3",x"13",x"13",x"ED",x"43",x"49",
x"5C",x"2A",x"5D",x"5C",x"EB",x"21",x"55",x"15",x"E5",x"2A",x"61",x"5C",x"37",x"ED",x"52",x"E5",
x"60",x"69",x"CD",x"6E",x"19",x"20",x"06",x"CD",x"B8",x"19",x"CD",x"E8",x"19",x"C1",x"79",x"3D",
x"B0",x"28",x"28",x"C5",x"03",x"03",x"03",x"03",x"2B",x"ED",x"5B",x"53",x"5C",x"D5",x"CD",x"55",
x"16",x"E1",x"22",x"53",x"5C",x"C1",x"C5",x"13",x"2A",x"61",x"5C",x"2B",x"2B",x"ED",x"B8",x"2A",
x"49",x"5C",x"EB",x"C1",x"70",x"2B",x"71",x"2B",x"73",x"2B",x"72",x"F1",x"C3",x"A2",x"12",x"F4",
x"09",x"A8",x"10",x"4B",x"F4",x"09",x"C4",x"15",x"53",x"81",x"0F",x"C4",x"15",x"52",x"F4",x"09",
x"C4",x"15",x"50",x"80",x"CF",x"12",x"01",x"00",x"06",x"00",x"0B",x"00",x"01",x"00",x"01",x"00",
x"06",x"00",x"10",x"00",x"FD",x"CB",x"02",x"6E",x"20",x"04",x"FD",x"CB",x"02",x"DE",x"CD",x"E6",
x"15",x"D8",x"28",x"FA",x"CF",x"07",x"D9",x"E5",x"2A",x"51",x"5C",x"23",x"23",x"18",x"08",x"1E",
x"30",x"83",x"D9",x"E5",x"2A",x"51",x"5C",x"5E",x"23",x"56",x"EB",x"CD",x"2C",x"16",x"E1",x"D9",
x"C9",x"87",x"C6",x"16",x"6F",x"26",x"5C",x"5E",x"23",x"56",x"7A",x"B3",x"20",x"02",x"CF",x"17",
x"1B",x"2A",x"4F",x"5C",x"19",x"22",x"51",x"5C",x"FD",x"CB",x"30",x"A6",x"23",x"23",x"23",x"23",
x"4E",x"21",x"2D",x"16",x"CD",x"DC",x"16",x"D0",x"16",x"00",x"5E",x"19",x"E9",x"4B",x"06",x"53",
x"12",x"50",x"1B",x"00",x"FD",x"CB",x"02",x"C6",x"FD",x"CB",x"01",x"AE",x"FD",x"CB",x"30",x"E6",
x"18",x"04",x"FD",x"CB",x"02",x"86",x"FD",x"CB",x"01",x"8E",x"C3",x"4D",x"0D",x"FD",x"CB",x"01",
x"CE",x"C9",x"01",x"01",x"00",x"E5",x"CD",x"05",x"1F",x"E1",x"CD",x"64",x"16",x"2A",x"65",x"5C",
x"EB",x"ED",x"B8",x"C9",x"F5",x"E5",x"21",x"4B",x"5C",x"3E",x"0E",x"5E",x"23",x"56",x"E3",x"A7",
x"ED",x"52",x"19",x"E3",x"30",x"09",x"D5",x"EB",x"09",x"EB",x"72",x"2B",x"73",x"23",x"D1",x"23",
x"3D",x"20",x"E8",x"EB",x"D1",x"F1",x"A7",x"ED",x"52",x"44",x"4D",x"03",x"19",x"EB",x"C9",x"00",
x"00",x"EB",x"11",x"8F",x"16",x"7E",x"E6",x"C0",x"20",x"F7",x"56",x"23",x"5E",x"C9",x"2A",x"63",
x"5C",x"2B",x"CD",x"55",x"16",x"23",x"23",x"C1",x"ED",x"43",x"61",x"5C",x"C1",x"EB",x"23",x"C9",
x"2A",x"59",x"5C",x"36",x"0D",x"22",x"5B",x"5C",x"23",x"36",x"80",x"23",x"22",x"61",x"5C",x"2A",
x"61",x"5C",x"22",x"63",x"5C",x"2A",x"63",x"5C",x"22",x"65",x"5C",x"E5",x"21",x"92",x"5C",x"22",
x"68",x"5C",x"E1",x"C9",x"ED",x"5B",x"59",x"5C",x"C3",x"E5",x"19",x"23",x"7E",x"A7",x"C8",x"B9",
x"23",x"20",x"F8",x"37",x"C9",x"CD",x"1E",x"17",x"CD",x"01",x"17",x"01",x"00",x"00",x"11",x"E2",
x"A3",x"EB",x"19",x"38",x"07",x"01",x"D4",x"15",x"09",x"4E",x"23",x"46",x"EB",x"71",x"23",x"70",
x"C9",x"E5",x"2A",x"4F",x"5C",x"09",x"23",x"23",x"23",x"4E",x"EB",x"21",x"16",x"17",x"CD",x"DC",
x"16",x"4E",x"06",x"00",x"09",x"E9",x"4B",x"05",x"53",x"03",x"50",x"01",x"E1",x"C9",x"CD",x"94",
x"1E",x"FE",x"10",x"38",x"02",x"CF",x"17",x"C6",x"03",x"07",x"21",x"10",x"5C",x"4F",x"06",x"00",
x"09",x"4E",x"23",x"46",x"2B",x"C9",x"EF",x"01",x"38",x"CD",x"1E",x"17",x"78",x"B1",x"28",x"16",
x"EB",x"2A",x"4F",x"5C",x"09",x"23",x"23",x"23",x"7E",x"EB",x"FE",x"4B",x"28",x"08",x"FE",x"53",
x"28",x"04",x"FE",x"50",x"20",x"CF",x"CD",x"5D",x"17",x"73",x"23",x"72",x"C9",x"E5",x"CD",x"F1",
x"2B",x"78",x"B1",x"20",x"02",x"CF",x"0E",x"C5",x"1A",x"E6",x"DF",x"4F",x"21",x"7A",x"17",x"CD",
x"DC",x"16",x"30",x"F1",x"4E",x"06",x"00",x"09",x"C1",x"E9",x"4B",x"06",x"53",x"08",x"50",x"0A",
x"00",x"1E",x"01",x"18",x"06",x"1E",x"06",x"18",x"02",x"1E",x"10",x"0B",x"78",x"B1",x"20",x"D5",
x"57",x"E1",x"C9",x"18",x"90",x"ED",x"73",x"3F",x"5C",x"FD",x"36",x"02",x"10",x"CD",x"AF",x"0D",
x"FD",x"CB",x"02",x"C6",x"FD",x"46",x"31",x"CD",x"44",x"0E",x"FD",x"CB",x"02",x"86",x"FD",x"CB",
x"30",x"C6",x"2A",x"49",x"5C",x"ED",x"5B",x"6C",x"5C",x"A7",x"ED",x"52",x"19",x"38",x"22",x"D5",
x"CD",x"6E",x"19",x"11",x"C0",x"02",x"EB",x"ED",x"52",x"E3",x"CD",x"6E",x"19",x"C1",x"C5",x"CD",
x"B8",x"19",x"C1",x"09",x"38",x"0E",x"EB",x"56",x"23",x"5E",x"2B",x"ED",x"53",x"6C",x"5C",x"18",
x"ED",x"22",x"6C",x"5C",x"2A",x"6C",x"5C",x"CD",x"6E",x"19",x"28",x"01",x"EB",x"CD",x"33",x"18",
x"FD",x"CB",x"02",x"A6",x"C9",x"3E",x"02",x"18",x"02",x"3E",x"02",x"FD",x"36",x"02",x"00",x"CD",
x"30",x"25",x"C4",x"01",x"16",x"DF",x"CD",x"70",x"20",x"38",x"14",x"DF",x"FE",x"3B",x"28",x"04",
x"FE",x"2C",x"20",x"06",x"E7",x"CD",x"82",x"1C",x"18",x"08",x"CD",x"E6",x"1C",x"18",x"03",x"CD",
x"DE",x"1C",x"CD",x"EE",x"1B",x"CD",x"99",x"1E",x"78",x"E6",x"3F",x"67",x"69",x"22",x"49",x"5C",
x"CD",x"6E",x"19",x"1E",x"01",x"CD",x"55",x"18",x"D7",x"FD",x"CB",x"02",x"66",x"28",x"F6",x"3A",
x"6B",x"5C",x"FD",x"96",x"4F",x"20",x"EE",x"AB",x"C8",x"E5",x"D5",x"21",x"6C",x"5C",x"CD",x"0F",
x"19",x"D1",x"E1",x"18",x"E0",x"ED",x"4B",x"49",x"5C",x"CD",x"80",x"19",x"16",x"3E",x"28",x"05",
x"11",x"00",x"00",x"CB",x"13",x"FD",x"73",x"2D",x"7E",x"FE",x"40",x"C1",x"D0",x"C5",x"CD",x"28",
x"1A",x"23",x"23",x"23",x"FD",x"CB",x"01",x"86",x"7A",x"A7",x"28",x"05",x"D7",x"FD",x"CB",x"01",
x"C6",x"D5",x"EB",x"FD",x"CB",x"30",x"96",x"21",x"3B",x"5C",x"CB",x"96",x"FD",x"CB",x"37",x"6E",
x"28",x"02",x"CB",x"D6",x"2A",x"5F",x"5C",x"A7",x"ED",x"52",x"20",x"05",x"3E",x"3F",x"CD",x"C1",
x"18",x"CD",x"E1",x"18",x"EB",x"7E",x"CD",x"B6",x"18",x"23",x"FE",x"0D",x"28",x"06",x"EB",x"CD",
x"37",x"19",x"18",x"E0",x"D1",x"C9",x"FE",x"0E",x"C0",x"23",x"23",x"23",x"23",x"23",x"23",x"7E",
x"C9",x"D9",x"2A",x"8F",x"5C",x"E5",x"CB",x"BC",x"CB",x"FD",x"22",x"8F",x"5C",x"21",x"91",x"5C",
x"56",x"D5",x"36",x"00",x"CD",x"F4",x"09",x"E1",x"FD",x"74",x"57",x"E1",x"22",x"8F",x"5C",x"D9",
x"C9",x"2A",x"5B",x"5C",x"A7",x"ED",x"52",x"C0",x"3A",x"41",x"5C",x"CB",x"07",x"28",x"04",x"C6",
x"43",x"18",x"16",x"21",x"3B",x"5C",x"CB",x"9E",x"3E",x"4B",x"CB",x"56",x"28",x"0B",x"CB",x"DE",
x"3C",x"FD",x"CB",x"30",x"5E",x"28",x"02",x"3E",x"43",x"D5",x"CD",x"C1",x"18",x"D1",x"C9",x"5E",
x"23",x"56",x"E5",x"EB",x"23",x"CD",x"6E",x"19",x"CD",x"95",x"16",x"E1",x"FD",x"CB",x"37",x"6E",
x"C0",x"72",x"2B",x"73",x"C9",x"7B",x"A7",x"F8",x"18",x"0D",x"AF",x"09",x"3C",x"38",x"FC",x"ED",
x"42",x"3D",x"28",x"F1",x"C3",x"EF",x"15",x"CD",x"1B",x"2D",x"30",x"30",x"FE",x"21",x"38",x"2C",
x"FD",x"CB",x"01",x"96",x"FE",x"CB",x"28",x"24",x"FE",x"3A",x"20",x"0E",x"FD",x"CB",x"37",x"6E",
x"20",x"16",x"FD",x"CB",x"30",x"56",x"28",x"14",x"18",x"0E",x"FE",x"22",x"20",x"0A",x"F5",x"3A",
x"6A",x"5C",x"EE",x"04",x"32",x"6A",x"5C",x"F1",x"FD",x"CB",x"01",x"D6",x"D7",x"C9",x"E5",x"2A",
x"53",x"5C",x"54",x"5D",x"C1",x"CD",x"80",x"19",x"D0",x"C5",x"CD",x"B8",x"19",x"EB",x"18",x"F4",
x"7E",x"B8",x"C0",x"23",x"7E",x"2B",x"B9",x"C9",x"23",x"23",x"23",x"22",x"5D",x"5C",x"0E",x"00",
x"15",x"C8",x"E7",x"BB",x"20",x"04",x"A7",x"C9",x"23",x"7E",x"CD",x"B6",x"18",x"22",x"5D",x"5C",
x"FE",x"22",x"20",x"01",x"0D",x"FE",x"3A",x"28",x"04",x"FE",x"CB",x"20",x"04",x"CB",x"41",x"28",
x"DF",x"FE",x"0D",x"20",x"E3",x"15",x"37",x"C9",x"E5",x"7E",x"FE",x"40",x"38",x"17",x"CB",x"6F",
x"28",x"14",x"87",x"FA",x"C7",x"19",x"3F",x"01",x"05",x"00",x"30",x"02",x"0E",x"12",x"17",x"23",
x"7E",x"30",x"FB",x"18",x"06",x"23",x"23",x"4E",x"23",x"46",x"23",x"09",x"D1",x"A7",x"ED",x"52",
x"44",x"4D",x"19",x"EB",x"C9",x"CD",x"DD",x"19",x"C5",x"78",x"2F",x"47",x"79",x"2F",x"4F",x"03",
x"CD",x"64",x"16",x"EB",x"E1",x"19",x"D5",x"ED",x"B0",x"E1",x"C9",x"2A",x"59",x"5C",x"2B",x"22",
x"5D",x"5C",x"E7",x"21",x"92",x"5C",x"22",x"65",x"5C",x"CD",x"3B",x"2D",x"CD",x"A2",x"2D",x"38",
x"04",x"21",x"F0",x"D8",x"09",x"DA",x"8A",x"1C",x"C3",x"C5",x"16",x"D5",x"E5",x"AF",x"CB",x"78",
x"20",x"20",x"60",x"69",x"1E",x"FF",x"18",x"08",x"D5",x"56",x"23",x"5E",x"E5",x"EB",x"1E",x"20",
x"01",x"18",x"FC",x"CD",x"2A",x"19",x"01",x"9C",x"FF",x"CD",x"2A",x"19",x"0E",x"F6",x"CD",x"2A",
x"19",x"7D",x"CD",x"EF",x"15",x"E1",x"D1",x"C9",x"B1",x"CB",x"BC",x"BF",x"C4",x"AF",x"B4",x"93",
x"91",x"92",x"95",x"98",x"98",x"98",x"98",x"98",x"98",x"98",x"7F",x"81",x"2E",x"6C",x"6E",x"70",
x"48",x"94",x"56",x"3F",x"41",x"2B",x"17",x"1F",x"37",x"77",x"44",x"0F",x"59",x"2B",x"43",x"2D",
x"51",x"3A",x"6D",x"42",x"0D",x"49",x"5C",x"44",x"15",x"5D",x"01",x"3D",x"02",x"06",x"00",x"67",
x"1E",x"06",x"CB",x"05",x"F0",x"1C",x"06",x"00",x"ED",x"1E",x"00",x"EE",x"1C",x"00",x"23",x"1F",
x"04",x"3D",x"06",x"CC",x"06",x"05",x"03",x"1D",x"04",x"00",x"AB",x"1D",x"05",x"CD",x"1F",x"05",
x"89",x"20",x"05",x"02",x"2C",x"05",x"B2",x"1B",x"00",x"B7",x"11",x"03",x"A1",x"1E",x"05",x"F9",
x"17",x"08",x"00",x"80",x"1E",x"03",x"4F",x"1E",x"00",x"5F",x"1E",x"03",x"AC",x"1E",x"00",x"6B",
x"0D",x"09",x"00",x"DC",x"22",x"06",x"00",x"3A",x"1F",x"05",x"ED",x"1D",x"05",x"27",x"1E",x"03",
x"42",x"1E",x"09",x"05",x"82",x"23",x"05",x"AC",x"0E",x"05",x"C9",x"1F",x"05",x"F5",x"17",x"0B",
x"0B",x"0B",x"0B",x"08",x"00",x"F8",x"03",x"09",x"05",x"20",x"23",x"07",x"07",x"07",x"07",x"07",
x"07",x"08",x"00",x"7A",x"1E",x"06",x"00",x"94",x"22",x"05",x"60",x"1F",x"06",x"2C",x"0A",x"00",
x"36",x"17",x"06",x"00",x"E5",x"16",x"0A",x"00",x"93",x"17",x"0A",x"2C",x"0A",x"00",x"93",x"17",
x"0A",x"00",x"93",x"17",x"00",x"93",x"17",x"FD",x"CB",x"01",x"BE",x"CD",x"FB",x"19",x"AF",x"32",
x"47",x"5C",x"3D",x"32",x"3A",x"5C",x"18",x"01",x"E7",x"CD",x"BF",x"16",x"FD",x"34",x"0D",x"FA",
x"8A",x"1C",x"DF",x"06",x"00",x"FE",x"0D",x"28",x"7A",x"FE",x"3A",x"28",x"EB",x"21",x"76",x"1B",
x"E5",x"4F",x"E7",x"79",x"D6",x"CE",x"DA",x"8A",x"1C",x"4F",x"21",x"48",x"1A",x"09",x"4E",x"09",
x"18",x"03",x"2A",x"74",x"5C",x"7E",x"23",x"22",x"74",x"5C",x"01",x"52",x"1B",x"C5",x"4F",x"FE",
x"20",x"30",x"0C",x"21",x"01",x"1C",x"06",x"00",x"09",x"4E",x"09",x"E5",x"DF",x"05",x"C9",x"DF",
x"B9",x"C2",x"8A",x"1C",x"E7",x"C9",x"CD",x"54",x"1F",x"38",x"02",x"CF",x"14",x"FD",x"CB",x"0A",
x"7E",x"20",x"71",x"2A",x"42",x"5C",x"CB",x"7C",x"28",x"14",x"21",x"FE",x"FF",x"22",x"45",x"5C",
x"2A",x"61",x"5C",x"2B",x"ED",x"5B",x"59",x"5C",x"1B",x"3A",x"44",x"5C",x"18",x"33",x"CD",x"6E",
x"19",x"3A",x"44",x"5C",x"28",x"19",x"A7",x"20",x"43",x"47",x"7E",x"E6",x"C0",x"78",x"28",x"0F",
x"CF",x"FF",x"C1",x"CD",x"30",x"25",x"C8",x"2A",x"55",x"5C",x"3E",x"C0",x"A6",x"C0",x"AF",x"FE",
x"01",x"CE",x"00",x"56",x"23",x"5E",x"ED",x"53",x"45",x"5C",x"23",x"5E",x"23",x"56",x"EB",x"19",
x"23",x"22",x"55",x"5C",x"EB",x"22",x"5D",x"5C",x"57",x"1E",x"00",x"FD",x"36",x"0A",x"FF",x"15",
x"FD",x"72",x"0D",x"CA",x"28",x"1B",x"14",x"CD",x"8B",x"19",x"28",x"08",x"CF",x"16",x"CD",x"30",
x"25",x"C0",x"C1",x"C1",x"DF",x"FE",x"0D",x"28",x"BA",x"FE",x"3A",x"CA",x"28",x"1B",x"C3",x"8A",
x"1C",x"0F",x"1D",x"4B",x"09",x"67",x"0B",x"7B",x"8E",x"71",x"B4",x"81",x"CF",x"CD",x"DE",x"1C",
x"BF",x"C1",x"CC",x"EE",x"1B",x"EB",x"2A",x"74",x"5C",x"4E",x"23",x"46",x"EB",x"C5",x"C9",x"CD",
x"B2",x"28",x"FD",x"36",x"37",x"00",x"30",x"08",x"FD",x"CB",x"37",x"CE",x"20",x"18",x"CF",x"01",
x"CC",x"96",x"29",x"FD",x"CB",x"01",x"76",x"20",x"0D",x"AF",x"CD",x"30",x"25",x"C4",x"F1",x"2B",
x"21",x"71",x"5C",x"B6",x"77",x"EB",x"ED",x"43",x"72",x"5C",x"22",x"4D",x"5C",x"C9",x"C1",x"CD",
x"56",x"1C",x"CD",x"EE",x"1B",x"C9",x"3A",x"3B",x"5C",x"F5",x"CD",x"FB",x"24",x"F1",x"FD",x"56",
x"01",x"AA",x"E6",x"40",x"20",x"24",x"CB",x"7A",x"C2",x"FF",x"2A",x"C9",x"CD",x"B2",x"28",x"F5",
x"79",x"F6",x"9F",x"3C",x"20",x"14",x"F1",x"18",x"A9",x"E7",x"CD",x"82",x"1C",x"FE",x"2C",x"20",
x"09",x"E7",x"CD",x"FB",x"24",x"FD",x"CB",x"01",x"76",x"C0",x"CF",x"0B",x"CD",x"FB",x"24",x"FD",
x"CB",x"01",x"76",x"C8",x"18",x"F4",x"FD",x"CB",x"01",x"7E",x"FD",x"CB",x"02",x"86",x"C4",x"4D",
x"0D",x"F1",x"3A",x"74",x"5C",x"D6",x"13",x"CD",x"FC",x"21",x"CD",x"EE",x"1B",x"2A",x"8F",x"5C",
x"22",x"8D",x"5C",x"21",x"91",x"5C",x"7E",x"07",x"AE",x"E6",x"AA",x"AE",x"77",x"C9",x"CD",x"30",
x"25",x"28",x"13",x"FD",x"CB",x"02",x"86",x"CD",x"4D",x"0D",x"21",x"90",x"5C",x"7E",x"F6",x"F8",
x"77",x"FD",x"CB",x"57",x"B6",x"DF",x"CD",x"E2",x"21",x"18",x"9F",x"C3",x"05",x"06",x"FE",x"0D",
x"28",x"04",x"FE",x"3A",x"20",x"9C",x"CD",x"30",x"25",x"C8",x"EF",x"A0",x"38",x"C9",x"CF",x"08",
x"C1",x"CD",x"30",x"25",x"28",x"0A",x"EF",x"02",x"38",x"EB",x"CD",x"E9",x"34",x"DA",x"B3",x"1B",
x"C3",x"29",x"1B",x"FE",x"CD",x"20",x"09",x"E7",x"CD",x"82",x"1C",x"CD",x"EE",x"1B",x"18",x"06",
x"CD",x"EE",x"1B",x"EF",x"A1",x"38",x"EF",x"C0",x"02",x"01",x"E0",x"01",x"38",x"CD",x"FF",x"2A",
x"22",x"68",x"5C",x"2B",x"7E",x"CB",x"FE",x"01",x"06",x"00",x"09",x"07",x"38",x"06",x"0E",x"0D",
x"CD",x"55",x"16",x"23",x"E5",x"EF",x"02",x"02",x"38",x"E1",x"EB",x"0E",x"0A",x"ED",x"B0",x"2A",
x"45",x"5C",x"EB",x"73",x"23",x"72",x"FD",x"56",x"0D",x"14",x"23",x"72",x"CD",x"DA",x"1D",x"D0",
x"FD",x"46",x"38",x"2A",x"45",x"5C",x"22",x"42",x"5C",x"3A",x"47",x"5C",x"ED",x"44",x"57",x"2A",
x"5D",x"5C",x"1E",x"F3",x"C5",x"ED",x"4B",x"55",x"5C",x"CD",x"86",x"1D",x"ED",x"43",x"55",x"5C",
x"C1",x"38",x"11",x"E7",x"F6",x"20",x"B8",x"28",x"03",x"E7",x"18",x"E8",x"E7",x"3E",x"01",x"92",
x"32",x"44",x"5C",x"C9",x"CF",x"11",x"7E",x"FE",x"3A",x"28",x"18",x"23",x"7E",x"E6",x"C0",x"37",
x"C0",x"46",x"23",x"4E",x"ED",x"43",x"42",x"5C",x"23",x"4E",x"23",x"46",x"E5",x"09",x"44",x"4D",
x"E1",x"16",x"00",x"C5",x"CD",x"8B",x"19",x"C1",x"D0",x"18",x"E0",x"FD",x"CB",x"37",x"4E",x"C2",
x"2E",x"1C",x"2A",x"4D",x"5C",x"CB",x"7E",x"28",x"1F",x"23",x"22",x"68",x"5C",x"EF",x"E0",x"E2",
x"0F",x"C0",x"02",x"38",x"CD",x"DA",x"1D",x"D8",x"2A",x"68",x"5C",x"11",x"0F",x"00",x"19",x"5E",
x"23",x"56",x"23",x"66",x"EB",x"C3",x"73",x"1E",x"CF",x"00",x"EF",x"E1",x"E0",x"E2",x"36",x"00",
x"02",x"01",x"03",x"37",x"00",x"04",x"38",x"A7",x"C9",x"38",x"37",x"C9",x"E7",x"CD",x"1F",x"1C",
x"CD",x"30",x"25",x"28",x"29",x"DF",x"22",x"5F",x"5C",x"2A",x"57",x"5C",x"7E",x"FE",x"2C",x"28",
x"09",x"1E",x"E4",x"CD",x"86",x"1D",x"30",x"02",x"CF",x"0D",x"CD",x"77",x"00",x"CD",x"56",x"1C",
x"DF",x"22",x"57",x"5C",x"2A",x"5F",x"5C",x"FD",x"36",x"26",x"00",x"CD",x"78",x"00",x"DF",x"FE",
x"2C",x"28",x"C9",x"CD",x"EE",x"1B",x"C9",x"CD",x"30",x"25",x"20",x"0B",x"CD",x"FB",x"24",x"FE",
x"2C",x"C4",x"EE",x"1B",x"E7",x"18",x"F5",x"3E",x"E4",x"47",x"ED",x"B9",x"11",x"00",x"02",x"C3",
x"8B",x"19",x"CD",x"99",x"1E",x"60",x"69",x"CD",x"6E",x"19",x"2B",x"22",x"57",x"5C",x"C9",x"CD",
x"99",x"1E",x"78",x"B1",x"20",x"04",x"ED",x"4B",x"78",x"5C",x"ED",x"43",x"76",x"5C",x"C9",x"2A",
x"6E",x"5C",x"FD",x"56",x"36",x"18",x"0C",x"CD",x"99",x"1E",x"60",x"69",x"16",x"00",x"7C",x"FE",
x"F0",x"30",x"2C",x"22",x"42",x"5C",x"FD",x"72",x"0A",x"C9",x"CD",x"85",x"1E",x"ED",x"79",x"C9",
x"CD",x"85",x"1E",x"02",x"C9",x"CD",x"D5",x"2D",x"38",x"15",x"28",x"02",x"ED",x"44",x"F5",x"CD",
x"99",x"1E",x"F1",x"C9",x"CD",x"D5",x"2D",x"18",x"03",x"CD",x"A2",x"2D",x"38",x"01",x"C8",x"CF",
x"0A",x"CD",x"67",x"1E",x"01",x"00",x"00",x"CD",x"45",x"1E",x"18",x"03",x"CD",x"99",x"1E",x"78",
x"B1",x"20",x"04",x"ED",x"4B",x"B2",x"5C",x"C5",x"ED",x"5B",x"4B",x"5C",x"2A",x"59",x"5C",x"2B",
x"CD",x"E5",x"19",x"CD",x"6B",x"0D",x"2A",x"65",x"5C",x"11",x"32",x"00",x"19",x"D1",x"ED",x"52",
x"30",x"08",x"2A",x"B4",x"5C",x"A7",x"ED",x"52",x"30",x"02",x"CF",x"15",x"EB",x"22",x"B2",x"5C",
x"D1",x"C1",x"36",x"3E",x"2B",x"F9",x"C5",x"ED",x"73",x"3D",x"5C",x"EB",x"E9",x"D1",x"FD",x"66",
x"0D",x"24",x"E3",x"33",x"ED",x"4B",x"45",x"5C",x"C5",x"E5",x"ED",x"73",x"3D",x"5C",x"D5",x"CD",
x"67",x"1E",x"01",x"14",x"00",x"2A",x"65",x"5C",x"09",x"38",x"0A",x"EB",x"21",x"50",x"00",x"19",
x"38",x"03",x"ED",x"72",x"D8",x"2E",x"03",x"C3",x"55",x"00",x"01",x"00",x"00",x"CD",x"05",x"1F",
x"44",x"4D",x"C9",x"C1",x"E1",x"D1",x"7A",x"FE",x"3E",x"28",x"0B",x"3B",x"E3",x"EB",x"ED",x"73",
x"3D",x"5C",x"C5",x"C3",x"73",x"1E",x"D5",x"E5",x"CF",x"06",x"CD",x"99",x"1E",x"76",x"0B",x"78",
x"B1",x"28",x"0C",x"78",x"A1",x"3C",x"20",x"01",x"03",x"FD",x"CB",x"01",x"6E",x"28",x"EE",x"FD",
x"CB",x"01",x"AE",x"C9",x"3E",x"7F",x"DB",x"FE",x"1F",x"D8",x"3E",x"FE",x"DB",x"FE",x"1F",x"C9",
x"CD",x"30",x"25",x"28",x"05",x"3E",x"CE",x"C3",x"39",x"1E",x"FD",x"CB",x"01",x"F6",x"CD",x"8D",
x"2C",x"30",x"16",x"E7",x"FE",x"24",x"20",x"05",x"FD",x"CB",x"01",x"B6",x"E7",x"FE",x"28",x"20",
x"3C",x"E7",x"FE",x"29",x"28",x"20",x"CD",x"8D",x"2C",x"D2",x"8A",x"1C",x"EB",x"E7",x"FE",x"24",
x"20",x"02",x"EB",x"E7",x"EB",x"01",x"06",x"00",x"CD",x"55",x"16",x"23",x"23",x"36",x"0E",x"FE",
x"2C",x"20",x"03",x"E7",x"18",x"E0",x"FE",x"29",x"20",x"13",x"E7",x"FE",x"3D",x"20",x"0E",x"E7",
x"3A",x"3B",x"5C",x"F5",x"CD",x"FB",x"24",x"F1",x"FD",x"AE",x"01",x"E6",x"40",x"C2",x"8A",x"1C",
x"CD",x"EE",x"1B",x"CD",x"30",x"25",x"E1",x"C8",x"E9",x"3E",x"02",x"18",x"02",x"3E",x"02",x"CD",
x"30",x"25",x"C4",x"01",x"16",x"CD",x"4D",x"0D",x"CD",x"DF",x"1F",x"CD",x"EE",x"1B",x"C9",x"DF",
x"CD",x"45",x"20",x"28",x"0D",x"CD",x"4E",x"20",x"28",x"FB",x"CD",x"FC",x"1F",x"CD",x"4E",x"20",
x"28",x"F3",x"FE",x"29",x"C8",x"CD",x"C3",x"1F",x"3E",x"0D",x"D7",x"C9",x"DF",x"FE",x"AC",x"20",
x"0D",x"CD",x"79",x"1C",x"CD",x"C3",x"1F",x"CD",x"07",x"23",x"3E",x"16",x"18",x"10",x"FE",x"AD",
x"20",x"12",x"E7",x"CD",x"82",x"1C",x"CD",x"C3",x"1F",x"CD",x"99",x"1E",x"3E",x"17",x"D7",x"79",
x"D7",x"78",x"D7",x"C9",x"CD",x"F2",x"21",x"D0",x"CD",x"70",x"20",x"D0",x"CD",x"FB",x"24",x"CD",
x"C3",x"1F",x"FD",x"CB",x"01",x"76",x"CC",x"F1",x"2B",x"C2",x"E3",x"2D",x"78",x"B1",x"0B",x"C8",
x"1A",x"13",x"D7",x"18",x"F7",x"FE",x"29",x"C8",x"FE",x"0D",x"C8",x"FE",x"3A",x"C9",x"DF",x"FE",
x"3B",x"28",x"14",x"FE",x"2C",x"20",x"0A",x"CD",x"30",x"25",x"28",x"0B",x"3E",x"06",x"D7",x"18",
x"06",x"FE",x"27",x"C0",x"CD",x"F5",x"1F",x"E7",x"CD",x"45",x"20",x"20",x"01",x"C1",x"BF",x"C9",
x"FE",x"23",x"37",x"C0",x"E7",x"CD",x"82",x"1C",x"A7",x"CD",x"C3",x"1F",x"CD",x"94",x"1E",x"FE",
x"10",x"D2",x"0E",x"16",x"CD",x"01",x"16",x"A7",x"C9",x"CD",x"30",x"25",x"28",x"08",x"3E",x"01",
x"CD",x"01",x"16",x"CD",x"6E",x"0D",x"FD",x"36",x"02",x"01",x"CD",x"C1",x"20",x"CD",x"EE",x"1B",
x"ED",x"4B",x"88",x"5C",x"3A",x"6B",x"5C",x"B8",x"38",x"03",x"0E",x"21",x"47",x"ED",x"43",x"88",
x"5C",x"3E",x"19",x"90",x"32",x"8C",x"5C",x"FD",x"CB",x"02",x"86",x"CD",x"D9",x"0D",x"C3",x"6E",
x"0D",x"CD",x"4E",x"20",x"28",x"FB",x"FE",x"28",x"20",x"0E",x"E7",x"CD",x"DF",x"1F",x"DF",x"FE",
x"29",x"C2",x"8A",x"1C",x"E7",x"C3",x"B2",x"21",x"FE",x"CA",x"20",x"11",x"E7",x"CD",x"1F",x"1C",
x"FD",x"CB",x"37",x"FE",x"FD",x"CB",x"01",x"76",x"C2",x"8A",x"1C",x"18",x"0D",x"CD",x"8D",x"2C",
x"D2",x"AF",x"21",x"CD",x"1F",x"1C",x"FD",x"CB",x"37",x"BE",x"CD",x"30",x"25",x"CA",x"B2",x"21",
x"CD",x"BF",x"16",x"21",x"71",x"5C",x"CB",x"B6",x"CB",x"EE",x"01",x"01",x"00",x"CB",x"7E",x"20",
x"0B",x"3A",x"3B",x"5C",x"E6",x"40",x"20",x"02",x"0E",x"03",x"B6",x"77",x"F7",x"36",x"0D",x"79",
x"0F",x"0F",x"30",x"05",x"3E",x"22",x"12",x"2B",x"77",x"22",x"5B",x"5C",x"FD",x"CB",x"37",x"7E",
x"20",x"2C",x"2A",x"5D",x"5C",x"E5",x"2A",x"3D",x"5C",x"E5",x"21",x"3A",x"21",x"E5",x"FD",x"CB",
x"30",x"66",x"28",x"04",x"ED",x"73",x"3D",x"5C",x"2A",x"61",x"5C",x"CD",x"A7",x"11",x"FD",x"36",
x"00",x"FF",x"CD",x"2C",x"0F",x"FD",x"CB",x"01",x"BE",x"CD",x"B9",x"21",x"18",x"03",x"CD",x"2C",
x"0F",x"FD",x"36",x"22",x"00",x"CD",x"D6",x"21",x"20",x"0A",x"CD",x"1D",x"11",x"ED",x"4B",x"82",
x"5C",x"CD",x"D9",x"0D",x"21",x"71",x"5C",x"CB",x"AE",x"CB",x"7E",x"CB",x"BE",x"20",x"1C",x"E1",
x"E1",x"22",x"3D",x"5C",x"E1",x"22",x"5F",x"5C",x"FD",x"CB",x"01",x"FE",x"CD",x"B9",x"21",x"2A",
x"5F",x"5C",x"FD",x"36",x"26",x"00",x"22",x"5D",x"5C",x"18",x"17",x"2A",x"63",x"5C",x"ED",x"5B",
x"61",x"5C",x"37",x"ED",x"52",x"44",x"4D",x"CD",x"B2",x"2A",x"CD",x"FF",x"2A",x"18",x"03",x"CD",
x"FC",x"1F",x"CD",x"4E",x"20",x"CA",x"C1",x"20",x"C9",x"2A",x"61",x"5C",x"22",x"5D",x"5C",x"DF",
x"FE",x"E2",x"28",x"0C",x"3A",x"71",x"5C",x"CD",x"59",x"1C",x"DF",x"FE",x"0D",x"C8",x"CF",x"0B",
x"CD",x"30",x"25",x"C8",x"CF",x"10",x"2A",x"51",x"5C",x"23",x"23",x"23",x"23",x"7E",x"FE",x"4B",
x"C9",x"E7",x"CD",x"F2",x"21",x"D8",x"DF",x"FE",x"2C",x"28",x"F6",x"FE",x"3B",x"28",x"F2",x"C3",
x"8A",x"1C",x"FE",x"D9",x"D8",x"FE",x"DF",x"3F",x"D8",x"F5",x"E7",x"F1",x"D6",x"C9",x"F5",x"CD",
x"82",x"1C",x"F1",x"A7",x"CD",x"C3",x"1F",x"F5",x"CD",x"94",x"1E",x"57",x"F1",x"D7",x"7A",x"D7",
x"C9",x"D6",x"11",x"CE",x"00",x"28",x"1D",x"D6",x"02",x"CE",x"00",x"28",x"56",x"FE",x"01",x"7A",
x"06",x"01",x"20",x"04",x"07",x"07",x"06",x"04",x"4F",x"7A",x"FE",x"02",x"30",x"16",x"79",x"21",
x"91",x"5C",x"18",x"38",x"7A",x"06",x"07",x"38",x"05",x"07",x"07",x"07",x"06",x"38",x"4F",x"7A",
x"FE",x"0A",x"38",x"02",x"CF",x"13",x"21",x"8F",x"5C",x"FE",x"08",x"38",x"0B",x"7E",x"28",x"07",
x"B0",x"2F",x"E6",x"24",x"28",x"01",x"78",x"4F",x"79",x"CD",x"6C",x"22",x"3E",x"07",x"BA",x"9F",
x"CD",x"6C",x"22",x"07",x"07",x"E6",x"50",x"47",x"3E",x"08",x"BA",x"9F",x"AE",x"A0",x"AE",x"77",
x"23",x"78",x"C9",x"9F",x"7A",x"0F",x"06",x"80",x"20",x"03",x"0F",x"06",x"40",x"4F",x"7A",x"FE",
x"08",x"28",x"04",x"FE",x"02",x"30",x"BD",x"79",x"21",x"8F",x"5C",x"CD",x"6C",x"22",x"79",x"0F",
x"0F",x"0F",x"18",x"D8",x"CD",x"94",x"1E",x"FE",x"08",x"30",x"A9",x"D3",x"FE",x"07",x"07",x"07",
x"CB",x"6F",x"20",x"02",x"EE",x"07",x"32",x"48",x"5C",x"C9",x"3E",x"AF",x"90",x"DA",x"F9",x"24",
x"47",x"A7",x"1F",x"37",x"1F",x"A7",x"1F",x"A8",x"E6",x"F8",x"A8",x"67",x"79",x"07",x"07",x"07",
x"A8",x"E6",x"C7",x"A8",x"07",x"07",x"6F",x"79",x"E6",x"07",x"C9",x"CD",x"07",x"23",x"CD",x"AA",
x"22",x"47",x"04",x"7E",x"07",x"10",x"FD",x"E6",x"01",x"C3",x"28",x"2D",x"CD",x"07",x"23",x"CD",
x"E5",x"22",x"C3",x"4D",x"0D",x"ED",x"43",x"7D",x"5C",x"CD",x"AA",x"22",x"47",x"04",x"3E",x"FE",
x"0F",x"10",x"FD",x"47",x"7E",x"FD",x"4E",x"57",x"CB",x"41",x"20",x"01",x"A0",x"CB",x"51",x"20",
x"02",x"A8",x"2F",x"77",x"C3",x"DB",x"0B",x"CD",x"14",x"23",x"47",x"C5",x"CD",x"14",x"23",x"59",
x"C1",x"51",x"4F",x"C9",x"CD",x"D5",x"2D",x"DA",x"F9",x"24",x"0E",x"01",x"C8",x"0E",x"FF",x"C9",
x"DF",x"FE",x"2C",x"C2",x"8A",x"1C",x"E7",x"CD",x"82",x"1C",x"CD",x"EE",x"1B",x"EF",x"2A",x"3D",
x"38",x"7E",x"FE",x"81",x"30",x"05",x"EF",x"02",x"38",x"18",x"A1",x"EF",x"A3",x"38",x"36",x"83",
x"EF",x"C5",x"02",x"38",x"CD",x"7D",x"24",x"C5",x"EF",x"31",x"E1",x"04",x"38",x"7E",x"FE",x"80",
x"30",x"08",x"EF",x"02",x"02",x"38",x"C1",x"C3",x"DC",x"22",x"EF",x"C2",x"01",x"C0",x"02",x"03",
x"01",x"E0",x"0F",x"C0",x"01",x"31",x"E0",x"01",x"31",x"E0",x"A0",x"C1",x"02",x"38",x"FD",x"34",
x"62",x"CD",x"94",x"1E",x"6F",x"E5",x"CD",x"94",x"1E",x"E1",x"67",x"22",x"7D",x"5C",x"C1",x"C3",
x"20",x"24",x"DF",x"FE",x"2C",x"28",x"06",x"CD",x"EE",x"1B",x"C3",x"77",x"24",x"E7",x"CD",x"82",
x"1C",x"CD",x"EE",x"1B",x"EF",x"C5",x"A2",x"04",x"1F",x"31",x"30",x"30",x"00",x"06",x"02",x"38",
x"C3",x"77",x"24",x"C0",x"02",x"C1",x"02",x"31",x"2A",x"E1",x"01",x"E1",x"2A",x"0F",x"E0",x"05",
x"2A",x"E0",x"01",x"3D",x"38",x"7E",x"FE",x"81",x"30",x"07",x"EF",x"02",x"02",x"38",x"C3",x"77",
x"24",x"CD",x"7D",x"24",x"C5",x"EF",x"02",x"E1",x"01",x"05",x"C1",x"02",x"01",x"31",x"E1",x"04",
x"C2",x"02",x"01",x"31",x"E1",x"04",x"E2",x"E5",x"E0",x"03",x"A2",x"04",x"31",x"1F",x"C5",x"02",
x"20",x"C0",x"02",x"C2",x"02",x"C1",x"E5",x"04",x"E0",x"E2",x"04",x"0F",x"E1",x"01",x"C1",x"02",
x"E0",x"04",x"E2",x"E5",x"04",x"03",x"C2",x"2A",x"E1",x"2A",x"0F",x"02",x"38",x"1A",x"FE",x"81",
x"C1",x"DA",x"77",x"24",x"C5",x"EF",x"01",x"38",x"3A",x"7D",x"5C",x"CD",x"28",x"2D",x"EF",x"C0",
x"0F",x"01",x"38",x"3A",x"7E",x"5C",x"CD",x"28",x"2D",x"EF",x"C5",x"0F",x"E0",x"E5",x"38",x"C1",
x"05",x"28",x"3C",x"18",x"14",x"EF",x"E1",x"31",x"E3",x"04",x"E2",x"E4",x"04",x"03",x"C1",x"02",
x"E4",x"04",x"E2",x"E3",x"04",x"0F",x"C2",x"02",x"38",x"C5",x"EF",x"C0",x"02",x"E1",x"0F",x"31",
x"38",x"3A",x"7D",x"5C",x"CD",x"28",x"2D",x"EF",x"03",x"E0",x"E2",x"0F",x"C0",x"01",x"E0",x"38",
x"3A",x"7E",x"5C",x"CD",x"28",x"2D",x"EF",x"03",x"38",x"CD",x"B7",x"24",x"C1",x"10",x"C6",x"EF",
x"02",x"02",x"01",x"38",x"3A",x"7D",x"5C",x"CD",x"28",x"2D",x"EF",x"03",x"01",x"38",x"3A",x"7E",
x"5C",x"CD",x"28",x"2D",x"EF",x"03",x"38",x"CD",x"B7",x"24",x"C3",x"4D",x"0D",x"EF",x"31",x"28",
x"34",x"32",x"00",x"01",x"05",x"E5",x"01",x"05",x"2A",x"38",x"CD",x"D5",x"2D",x"38",x"06",x"E6",
x"FC",x"C6",x"04",x"30",x"02",x"3E",x"FC",x"F5",x"CD",x"28",x"2D",x"EF",x"E5",x"01",x"05",x"31",
x"1F",x"C4",x"02",x"31",x"A2",x"04",x"1F",x"C1",x"01",x"C0",x"02",x"31",x"04",x"31",x"0F",x"A1",
x"03",x"1B",x"C3",x"02",x"38",x"C1",x"C9",x"CD",x"07",x"23",x"79",x"B8",x"30",x"06",x"69",x"D5",
x"AF",x"5F",x"18",x"07",x"B1",x"C8",x"68",x"41",x"D5",x"16",x"00",x"60",x"78",x"1F",x"85",x"38",
x"03",x"BC",x"38",x"07",x"94",x"4F",x"D9",x"C1",x"C5",x"18",x"04",x"4F",x"D5",x"D9",x"C1",x"2A",
x"7D",x"5C",x"78",x"84",x"47",x"79",x"3C",x"85",x"38",x"0D",x"28",x"0D",x"3D",x"4F",x"CD",x"E5",
x"22",x"D9",x"79",x"10",x"D9",x"D1",x"C9",x"28",x"F3",x"CF",x"0A",x"DF",x"06",x"00",x"C5",x"4F",
x"21",x"96",x"25",x"CD",x"DC",x"16",x"79",x"D2",x"84",x"26",x"06",x"00",x"4E",x"09",x"E9",x"CD",
x"74",x"00",x"03",x"FE",x"0D",x"CA",x"8A",x"1C",x"FE",x"22",x"20",x"F3",x"CD",x"74",x"00",x"FE",
x"22",x"C9",x"E7",x"FE",x"28",x"20",x"06",x"CD",x"79",x"1C",x"DF",x"FE",x"29",x"C2",x"8A",x"1C",
x"FD",x"CB",x"01",x"7E",x"C9",x"CD",x"07",x"23",x"2A",x"36",x"5C",x"11",x"00",x"01",x"19",x"79",
x"0F",x"0F",x"0F",x"E6",x"E0",x"A8",x"5F",x"79",x"E6",x"18",x"EE",x"40",x"57",x"06",x"60",x"C5",
x"D5",x"E5",x"1A",x"AE",x"28",x"04",x"3C",x"20",x"1A",x"3D",x"4F",x"06",x"07",x"14",x"23",x"1A",
x"AE",x"A9",x"20",x"0F",x"10",x"F7",x"C1",x"C1",x"C1",x"3E",x"80",x"90",x"01",x"01",x"00",x"F7",
x"12",x"18",x"0A",x"E1",x"11",x"08",x"00",x"19",x"D1",x"C1",x"10",x"D3",x"48",x"C3",x"B2",x"2A",
x"CD",x"07",x"23",x"79",x"0F",x"0F",x"0F",x"4F",x"E6",x"E0",x"A8",x"6F",x"79",x"E6",x"03",x"EE",
x"58",x"67",x"7E",x"C3",x"28",x"2D",x"22",x"1C",x"28",x"4F",x"2E",x"F2",x"2B",x"12",x"A8",x"56",
x"A5",x"57",x"A7",x"84",x"A6",x"8F",x"C4",x"E6",x"AA",x"BF",x"AB",x"C7",x"A9",x"CE",x"00",x"E7",
x"C3",x"FF",x"24",x"DF",x"23",x"E5",x"01",x"00",x"00",x"CD",x"0F",x"25",x"20",x"1B",x"CD",x"0F",
x"25",x"28",x"FB",x"CD",x"30",x"25",x"28",x"11",x"F7",x"E1",x"D5",x"7E",x"23",x"12",x"13",x"FE",
x"22",x"20",x"F8",x"7E",x"23",x"FE",x"22",x"28",x"F2",x"0B",x"D1",x"21",x"3B",x"5C",x"CB",x"B6",
x"CB",x"7E",x"C4",x"B2",x"2A",x"C3",x"12",x"27",x"E7",x"CD",x"FB",x"24",x"FE",x"29",x"C2",x"8A",
x"1C",x"E7",x"C3",x"12",x"27",x"C3",x"BD",x"27",x"CD",x"30",x"25",x"28",x"28",x"ED",x"4B",x"76",
x"5C",x"CD",x"2B",x"2D",x"EF",x"A1",x"0F",x"34",x"37",x"16",x"04",x"34",x"80",x"41",x"00",x"00",
x"80",x"32",x"02",x"A1",x"03",x"31",x"38",x"CD",x"A2",x"2D",x"ED",x"43",x"76",x"5C",x"7E",x"A7",
x"28",x"03",x"D6",x"10",x"77",x"18",x"09",x"CD",x"30",x"25",x"28",x"04",x"EF",x"A3",x"38",x"34",
x"E7",x"C3",x"C3",x"26",x"01",x"5A",x"10",x"E7",x"FE",x"23",x"CA",x"0D",x"27",x"21",x"3B",x"5C",
x"CB",x"B6",x"CB",x"7E",x"28",x"1F",x"CD",x"8E",x"02",x"0E",x"00",x"20",x"13",x"CD",x"1E",x"03",
x"30",x"0E",x"15",x"5F",x"CD",x"33",x"03",x"F5",x"01",x"01",x"00",x"F7",x"F1",x"12",x"0E",x"01",
x"06",x"00",x"CD",x"B2",x"2A",x"C3",x"12",x"27",x"CD",x"22",x"25",x"C4",x"35",x"25",x"E7",x"C3",
x"DB",x"25",x"CD",x"22",x"25",x"C4",x"80",x"25",x"E7",x"18",x"48",x"CD",x"22",x"25",x"C4",x"CB",
x"22",x"E7",x"18",x"3F",x"CD",x"88",x"2C",x"30",x"56",x"FE",x"41",x"30",x"3C",x"CD",x"30",x"25",
x"20",x"23",x"CD",x"9B",x"2C",x"DF",x"01",x"06",x"00",x"CD",x"55",x"16",x"23",x"36",x"0E",x"23",
x"EB",x"2A",x"65",x"5C",x"0E",x"05",x"A7",x"ED",x"42",x"22",x"65",x"5C",x"ED",x"B0",x"EB",x"2B",
x"CD",x"77",x"00",x"18",x"0E",x"DF",x"23",x"7E",x"FE",x"0E",x"20",x"FA",x"23",x"CD",x"B4",x"33",
x"22",x"5D",x"5C",x"FD",x"CB",x"01",x"F6",x"18",x"14",x"CD",x"B2",x"28",x"DA",x"2E",x"1C",x"CC",
x"96",x"29",x"3A",x"3B",x"5C",x"FE",x"C0",x"38",x"04",x"23",x"CD",x"B4",x"33",x"18",x"33",x"01",
x"DB",x"09",x"FE",x"2D",x"28",x"27",x"01",x"18",x"10",x"FE",x"AE",x"28",x"20",x"D6",x"AF",x"DA",
x"8A",x"1C",x"01",x"F0",x"04",x"FE",x"14",x"28",x"14",x"D2",x"8A",x"1C",x"06",x"10",x"C6",x"DC",
x"4F",x"FE",x"DF",x"30",x"02",x"CB",x"B1",x"FE",x"EE",x"38",x"02",x"CB",x"B9",x"C5",x"E7",x"C3",
x"FF",x"24",x"DF",x"FE",x"28",x"20",x"0C",x"FD",x"CB",x"01",x"76",x"20",x"17",x"CD",x"52",x"2A",
x"E7",x"18",x"F0",x"06",x"00",x"4F",x"21",x"95",x"27",x"CD",x"DC",x"16",x"30",x"06",x"4E",x"21",
x"ED",x"26",x"09",x"46",x"D1",x"7A",x"B8",x"38",x"3A",x"A7",x"CA",x"18",x"00",x"C5",x"21",x"3B",
x"5C",x"7B",x"FE",x"ED",x"20",x"06",x"CB",x"76",x"20",x"02",x"1E",x"99",x"D5",x"CD",x"30",x"25",
x"28",x"09",x"7B",x"E6",x"3F",x"47",x"EF",x"3B",x"38",x"18",x"09",x"7B",x"FD",x"AE",x"01",x"E6",
x"40",x"C2",x"8A",x"1C",x"D1",x"21",x"3B",x"5C",x"CB",x"F6",x"CB",x"7B",x"20",x"02",x"CB",x"B6",
x"C1",x"18",x"C1",x"D5",x"79",x"FD",x"CB",x"01",x"76",x"20",x"15",x"E6",x"3F",x"C6",x"08",x"4F",
x"FE",x"10",x"20",x"04",x"CB",x"F1",x"18",x"08",x"38",x"D7",x"FE",x"17",x"28",x"02",x"CB",x"F9",
x"C5",x"E7",x"C3",x"FF",x"24",x"2B",x"CF",x"2D",x"C3",x"2A",x"C4",x"2F",x"C5",x"5E",x"C6",x"3D",
x"CE",x"3E",x"CC",x"3C",x"CD",x"C7",x"C9",x"C8",x"CA",x"C9",x"CB",x"C5",x"C7",x"C6",x"C8",x"00",
x"06",x"08",x"08",x"0A",x"02",x"03",x"05",x"05",x"05",x"05",x"05",x"05",x"06",x"CD",x"30",x"25",
x"20",x"35",x"E7",x"CD",x"8D",x"2C",x"D2",x"8A",x"1C",x"E7",x"FE",x"24",x"F5",x"20",x"01",x"E7",
x"FE",x"28",x"20",x"12",x"E7",x"FE",x"29",x"28",x"10",x"CD",x"FB",x"24",x"DF",x"FE",x"2C",x"20",
x"03",x"E7",x"18",x"F5",x"FE",x"29",x"C2",x"8A",x"1C",x"E7",x"21",x"3B",x"5C",x"CB",x"B6",x"F1",
x"28",x"02",x"CB",x"F6",x"C3",x"12",x"27",x"E7",x"E6",x"DF",x"47",x"E7",x"D6",x"24",x"4F",x"20",
x"01",x"E7",x"E7",x"E5",x"2A",x"53",x"5C",x"2B",x"11",x"CE",x"00",x"C5",x"CD",x"86",x"1D",x"C1",
x"30",x"02",x"CF",x"18",x"E5",x"CD",x"AB",x"28",x"E6",x"DF",x"B8",x"20",x"08",x"CD",x"AB",x"28",
x"D6",x"24",x"B9",x"28",x"0C",x"E1",x"2B",x"11",x"00",x"02",x"C5",x"CD",x"8B",x"19",x"C1",x"18",
x"D7",x"A7",x"CC",x"AB",x"28",x"D1",x"D1",x"ED",x"53",x"5D",x"5C",x"CD",x"AB",x"28",x"E5",x"FE",
x"29",x"28",x"42",x"23",x"7E",x"FE",x"0E",x"16",x"40",x"28",x"07",x"2B",x"CD",x"AB",x"28",x"23",
x"16",x"00",x"23",x"E5",x"D5",x"CD",x"FB",x"24",x"F1",x"FD",x"AE",x"01",x"E6",x"40",x"20",x"2B",
x"E1",x"EB",x"2A",x"65",x"5C",x"01",x"05",x"00",x"ED",x"42",x"22",x"65",x"5C",x"ED",x"B0",x"EB",
x"2B",x"CD",x"AB",x"28",x"FE",x"29",x"28",x"0D",x"E5",x"DF",x"FE",x"2C",x"20",x"0D",x"E7",x"E1",
x"CD",x"AB",x"28",x"18",x"BE",x"E5",x"DF",x"FE",x"29",x"28",x"02",x"CF",x"19",x"D1",x"EB",x"22",
x"5D",x"5C",x"2A",x"0B",x"5C",x"E3",x"22",x"0B",x"5C",x"D5",x"E7",x"E7",x"CD",x"FB",x"24",x"E1",
x"22",x"5D",x"5C",x"E1",x"22",x"0B",x"5C",x"E7",x"C3",x"12",x"27",x"23",x"7E",x"FE",x"21",x"38",
x"FA",x"C9",x"FD",x"CB",x"01",x"F6",x"DF",x"CD",x"8D",x"2C",x"D2",x"8A",x"1C",x"E5",x"E6",x"1F",
x"4F",x"E7",x"E5",x"FE",x"28",x"28",x"28",x"CB",x"F1",x"FE",x"24",x"28",x"11",x"CB",x"E9",x"CD",
x"88",x"2C",x"30",x"0F",x"CD",x"88",x"2C",x"30",x"16",x"CB",x"B1",x"E7",x"18",x"F6",x"E7",x"FD",
x"CB",x"01",x"B6",x"3A",x"0C",x"5C",x"A7",x"28",x"06",x"CD",x"30",x"25",x"C2",x"51",x"29",x"41",
x"CD",x"30",x"25",x"20",x"08",x"79",x"E6",x"E0",x"CB",x"FF",x"4F",x"18",x"37",x"2A",x"4B",x"5C",
x"7E",x"E6",x"7F",x"28",x"2D",x"B9",x"20",x"22",x"17",x"87",x"F2",x"3F",x"29",x"38",x"30",x"D1",
x"D5",x"E5",x"23",x"1A",x"13",x"FE",x"20",x"28",x"FA",x"F6",x"20",x"BE",x"28",x"F4",x"F6",x"80",
x"BE",x"20",x"06",x"1A",x"CD",x"88",x"2C",x"30",x"15",x"E1",x"C5",x"CD",x"B8",x"19",x"EB",x"C1",
x"18",x"CE",x"CB",x"F8",x"D1",x"DF",x"FE",x"28",x"28",x"09",x"CB",x"E8",x"18",x"0D",x"D1",x"D1",
x"D1",x"E5",x"DF",x"CD",x"88",x"2C",x"30",x"03",x"E7",x"18",x"F8",x"E1",x"CB",x"10",x"CB",x"70",
x"C9",x"2A",x"0B",x"5C",x"7E",x"FE",x"29",x"CA",x"EF",x"28",x"7E",x"F6",x"60",x"47",x"23",x"7E",
x"FE",x"0E",x"28",x"07",x"2B",x"CD",x"AB",x"28",x"23",x"CB",x"A8",x"78",x"B9",x"28",x"12",x"23",
x"23",x"23",x"23",x"23",x"CD",x"AB",x"28",x"FE",x"29",x"CA",x"EF",x"28",x"CD",x"AB",x"28",x"18",
x"D9",x"CB",x"69",x"20",x"0C",x"23",x"ED",x"5B",x"65",x"5C",x"CD",x"C0",x"33",x"EB",x"22",x"65",
x"5C",x"D1",x"D1",x"AF",x"3C",x"C9",x"AF",x"47",x"CB",x"79",x"20",x"4B",x"CB",x"7E",x"20",x"0E",
x"3C",x"23",x"4E",x"23",x"46",x"23",x"EB",x"CD",x"B2",x"2A",x"DF",x"C3",x"49",x"2A",x"23",x"23",
x"23",x"46",x"CB",x"71",x"28",x"0A",x"05",x"28",x"E8",x"EB",x"DF",x"FE",x"28",x"20",x"61",x"EB",
x"EB",x"18",x"24",x"E5",x"DF",x"E1",x"FE",x"2C",x"28",x"20",x"CB",x"79",x"28",x"52",x"CB",x"71",
x"20",x"06",x"FE",x"29",x"20",x"3C",x"E7",x"C9",x"FE",x"29",x"28",x"6C",x"FE",x"CC",x"20",x"32",
x"DF",x"2B",x"22",x"5D",x"5C",x"18",x"5E",x"21",x"00",x"00",x"E5",x"E7",x"E1",x"79",x"FE",x"C0",
x"20",x"09",x"DF",x"FE",x"29",x"28",x"51",x"FE",x"CC",x"28",x"E5",x"C5",x"E5",x"CD",x"EE",x"2A",
x"E3",x"EB",x"CD",x"CC",x"2A",x"38",x"19",x"0B",x"CD",x"F4",x"2A",x"09",x"D1",x"C1",x"10",x"B3",
x"CB",x"79",x"20",x"66",x"E5",x"CB",x"71",x"20",x"13",x"42",x"4B",x"DF",x"FE",x"29",x"28",x"02",
x"CF",x"02",x"E7",x"E1",x"11",x"05",x"00",x"CD",x"F4",x"2A",x"09",x"C9",x"CD",x"EE",x"2A",x"E3",
x"CD",x"F4",x"2A",x"C1",x"09",x"23",x"42",x"4B",x"EB",x"CD",x"B1",x"2A",x"DF",x"FE",x"29",x"28",
x"07",x"FE",x"2C",x"20",x"DB",x"CD",x"52",x"2A",x"E7",x"FE",x"28",x"28",x"F8",x"FD",x"CB",x"01",
x"B6",x"C9",x"CD",x"30",x"25",x"C4",x"F1",x"2B",x"E7",x"FE",x"29",x"28",x"50",x"D5",x"AF",x"F5",
x"C5",x"11",x"01",x"00",x"DF",x"E1",x"FE",x"CC",x"28",x"17",x"F1",x"CD",x"CD",x"2A",x"F5",x"50",
x"59",x"E5",x"DF",x"E1",x"FE",x"CC",x"28",x"09",x"FE",x"29",x"C2",x"8A",x"1C",x"62",x"6B",x"18",
x"13",x"E5",x"E7",x"E1",x"FE",x"29",x"28",x"0C",x"F1",x"CD",x"CD",x"2A",x"F5",x"DF",x"60",x"69",
x"FE",x"29",x"20",x"E6",x"F1",x"E3",x"19",x"2B",x"E3",x"A7",x"ED",x"52",x"01",x"00",x"00",x"38",
x"07",x"23",x"A7",x"FA",x"20",x"2A",x"44",x"4D",x"D1",x"FD",x"CB",x"01",x"B6",x"CD",x"30",x"25",
x"C8",x"AF",x"FD",x"CB",x"01",x"B6",x"C5",x"CD",x"A9",x"33",x"C1",x"2A",x"65",x"5C",x"77",x"23",
x"73",x"23",x"72",x"23",x"71",x"23",x"70",x"23",x"22",x"65",x"5C",x"C9",x"AF",x"D5",x"E5",x"F5",
x"CD",x"82",x"1C",x"F1",x"CD",x"30",x"25",x"28",x"12",x"F5",x"CD",x"99",x"1E",x"D1",x"78",x"B1",
x"37",x"28",x"05",x"E1",x"E5",x"A7",x"ED",x"42",x"7A",x"DE",x"00",x"E1",x"D1",x"C9",x"EB",x"23",
x"5E",x"23",x"56",x"C9",x"CD",x"30",x"25",x"C8",x"CD",x"A9",x"30",x"DA",x"15",x"1F",x"C9",x"2A",
x"4D",x"5C",x"FD",x"CB",x"37",x"4E",x"28",x"5E",x"01",x"05",x"00",x"03",x"23",x"7E",x"FE",x"20",
x"28",x"FA",x"30",x"0B",x"FE",x"10",x"38",x"11",x"FE",x"16",x"30",x"0D",x"23",x"18",x"ED",x"CD",
x"88",x"2C",x"38",x"E7",x"FE",x"24",x"CA",x"C0",x"2B",x"79",x"2A",x"59",x"5C",x"2B",x"CD",x"55",
x"16",x"23",x"23",x"EB",x"D5",x"2A",x"4D",x"5C",x"1B",x"D6",x"06",x"47",x"28",x"11",x"23",x"7E",
x"FE",x"21",x"38",x"FA",x"F6",x"20",x"13",x"12",x"10",x"F4",x"F6",x"80",x"12",x"3E",x"C0",x"2A",
x"4D",x"5C",x"AE",x"F6",x"20",x"E1",x"CD",x"EA",x"2B",x"E5",x"EF",x"02",x"38",x"E1",x"01",x"05",
x"00",x"A7",x"ED",x"42",x"18",x"40",x"FD",x"CB",x"01",x"76",x"28",x"06",x"11",x"06",x"00",x"19",
x"18",x"E7",x"2A",x"4D",x"5C",x"ED",x"4B",x"72",x"5C",x"FD",x"CB",x"37",x"46",x"20",x"30",x"78",
x"B1",x"C8",x"E5",x"F7",x"D5",x"C5",x"54",x"5D",x"23",x"36",x"20",x"ED",x"B8",x"E5",x"CD",x"F1",
x"2B",x"E1",x"E3",x"A7",x"ED",x"42",x"09",x"30",x"02",x"44",x"4D",x"E3",x"EB",x"78",x"B1",x"28",
x"02",x"ED",x"B0",x"C1",x"D1",x"E1",x"EB",x"78",x"B1",x"C8",x"D5",x"ED",x"B0",x"E1",x"C9",x"2B",
x"2B",x"2B",x"7E",x"E5",x"C5",x"CD",x"C6",x"2B",x"C1",x"E1",x"03",x"03",x"03",x"C3",x"E8",x"19",
x"3E",x"DF",x"2A",x"4D",x"5C",x"A6",x"F5",x"CD",x"F1",x"2B",x"EB",x"09",x"C5",x"2B",x"22",x"4D",
x"5C",x"03",x"03",x"03",x"2A",x"59",x"5C",x"2B",x"CD",x"55",x"16",x"2A",x"4D",x"5C",x"C1",x"C5",
x"03",x"ED",x"B8",x"EB",x"23",x"C1",x"70",x"2B",x"71",x"F1",x"2B",x"77",x"2A",x"59",x"5C",x"2B",
x"C9",x"2A",x"65",x"5C",x"2B",x"46",x"2B",x"4E",x"2B",x"56",x"2B",x"5E",x"2B",x"7E",x"22",x"65",
x"5C",x"C9",x"CD",x"B2",x"28",x"C2",x"8A",x"1C",x"CD",x"30",x"25",x"20",x"08",x"CB",x"B1",x"CD",
x"96",x"29",x"CD",x"EE",x"1B",x"38",x"08",x"C5",x"CD",x"B8",x"19",x"CD",x"E8",x"19",x"C1",x"CB",
x"F9",x"06",x"00",x"C5",x"21",x"01",x"00",x"CB",x"71",x"20",x"02",x"2E",x"05",x"EB",x"E7",x"26",
x"FF",x"CD",x"CC",x"2A",x"DA",x"20",x"2A",x"E1",x"C5",x"24",x"E5",x"60",x"69",x"CD",x"F4",x"2A",
x"EB",x"DF",x"FE",x"2C",x"28",x"E8",x"FE",x"29",x"20",x"BB",x"E7",x"C1",x"79",x"68",x"26",x"00",
x"23",x"23",x"29",x"19",x"DA",x"15",x"1F",x"D5",x"C5",x"E5",x"44",x"4D",x"2A",x"59",x"5C",x"2B",
x"CD",x"55",x"16",x"23",x"77",x"C1",x"0B",x"0B",x"0B",x"23",x"71",x"23",x"70",x"C1",x"78",x"23",
x"77",x"62",x"6B",x"1B",x"36",x"00",x"CB",x"71",x"28",x"02",x"36",x"20",x"C1",x"ED",x"B8",x"C1",
x"70",x"2B",x"71",x"2B",x"3D",x"20",x"F8",x"C9",x"CD",x"1B",x"2D",x"3F",x"D8",x"FE",x"41",x"3F",
x"D0",x"FE",x"5B",x"D8",x"FE",x"61",x"3F",x"D0",x"FE",x"7B",x"C9",x"FE",x"C4",x"20",x"19",x"11",
x"00",x"00",x"E7",x"D6",x"31",x"CE",x"00",x"20",x"0A",x"EB",x"3F",x"ED",x"6A",x"DA",x"AD",x"31",
x"EB",x"18",x"EF",x"42",x"4B",x"C3",x"2B",x"2D",x"FE",x"2E",x"28",x"0F",x"CD",x"3B",x"2D",x"FE",
x"2E",x"20",x"28",x"E7",x"CD",x"1B",x"2D",x"38",x"22",x"18",x"0A",x"E7",x"CD",x"1B",x"2D",x"DA",
x"8A",x"1C",x"EF",x"A0",x"38",x"EF",x"A1",x"C0",x"02",x"38",x"DF",x"CD",x"22",x"2D",x"38",x"0B",
x"EF",x"E0",x"A4",x"05",x"C0",x"04",x"0F",x"38",x"E7",x"18",x"EF",x"FE",x"45",x"28",x"03",x"FE",
x"65",x"C0",x"06",x"FF",x"E7",x"FE",x"2B",x"28",x"05",x"FE",x"2D",x"20",x"02",x"04",x"E7",x"CD",
x"1B",x"2D",x"38",x"CB",x"C5",x"CD",x"3B",x"2D",x"CD",x"D5",x"2D",x"C1",x"DA",x"AD",x"31",x"A7",
x"FA",x"AD",x"31",x"04",x"28",x"02",x"ED",x"44",x"C3",x"4F",x"2D",x"FE",x"30",x"D8",x"FE",x"3A",
x"3F",x"C9",x"CD",x"1B",x"2D",x"D8",x"D6",x"30",x"4F",x"06",x"00",x"FD",x"21",x"3A",x"5C",x"AF",
x"5F",x"51",x"48",x"47",x"CD",x"B6",x"2A",x"EF",x"38",x"A7",x"C9",x"F5",x"EF",x"A0",x"38",x"F1",
x"CD",x"22",x"2D",x"D8",x"EF",x"01",x"A4",x"04",x"0F",x"38",x"CD",x"74",x"00",x"18",x"F1",x"07",
x"0F",x"30",x"02",x"2F",x"3C",x"F5",x"21",x"92",x"5C",x"CD",x"0B",x"35",x"EF",x"A4",x"38",x"F1",
x"CB",x"3F",x"30",x"0D",x"F5",x"EF",x"C1",x"E0",x"00",x"04",x"04",x"33",x"02",x"05",x"E1",x"38",
x"F1",x"28",x"08",x"F5",x"EF",x"31",x"04",x"38",x"F1",x"18",x"E5",x"EF",x"02",x"38",x"C9",x"23",
x"4E",x"23",x"7E",x"A9",x"91",x"5F",x"23",x"7E",x"89",x"A9",x"57",x"C9",x"0E",x"00",x"E5",x"36",
x"00",x"23",x"71",x"23",x"7B",x"A9",x"91",x"77",x"23",x"7A",x"89",x"A9",x"77",x"23",x"36",x"00",
x"E1",x"C9",x"EF",x"38",x"7E",x"A7",x"28",x"05",x"EF",x"A2",x"0F",x"27",x"38",x"EF",x"02",x"38",
x"E5",x"D5",x"EB",x"46",x"CD",x"7F",x"2D",x"AF",x"90",x"CB",x"79",x"42",x"4B",x"7B",x"D1",x"E1",
x"C9",x"57",x"17",x"9F",x"5F",x"4F",x"AF",x"47",x"CD",x"B6",x"2A",x"EF",x"34",x"EF",x"1A",x"20",
x"9A",x"85",x"04",x"27",x"38",x"CD",x"A2",x"2D",x"D8",x"F5",x"05",x"04",x"28",x"03",x"F1",x"37",
x"C9",x"F1",x"C9",x"EF",x"31",x"36",x"00",x"0B",x"31",x"37",x"00",x"0D",x"02",x"38",x"3E",x"30",
x"D7",x"C9",x"2A",x"38",x"3E",x"2D",x"D7",x"EF",x"A0",x"C3",x"C4",x"C5",x"02",x"38",x"D9",x"E5",
x"D9",x"EF",x"31",x"27",x"C2",x"03",x"E2",x"01",x"C2",x"02",x"38",x"7E",x"A7",x"20",x"47",x"CD",
x"7F",x"2D",x"06",x"10",x"7A",x"A7",x"20",x"06",x"B3",x"28",x"09",x"53",x"06",x"08",x"D5",x"D9",
x"D1",x"D9",x"18",x"57",x"EF",x"E2",x"38",x"7E",x"D6",x"7E",x"CD",x"C1",x"2D",x"57",x"3A",x"AC",
x"5C",x"92",x"32",x"AC",x"5C",x"7A",x"CD",x"4F",x"2D",x"EF",x"31",x"27",x"C1",x"03",x"E1",x"38",
x"CD",x"D5",x"2D",x"E5",x"32",x"A1",x"5C",x"3D",x"17",x"9F",x"3C",x"21",x"AB",x"5C",x"77",x"23",
x"86",x"77",x"E1",x"C3",x"CF",x"2E",x"D6",x"80",x"FE",x"1C",x"38",x"13",x"CD",x"C1",x"2D",x"D6",
x"07",x"47",x"21",x"AC",x"5C",x"86",x"77",x"78",x"ED",x"44",x"CD",x"4F",x"2D",x"18",x"92",x"EB",
x"CD",x"BA",x"2F",x"D9",x"CB",x"FA",x"7D",x"D9",x"D6",x"80",x"47",x"CB",x"23",x"CB",x"12",x"D9",
x"CB",x"13",x"CB",x"12",x"D9",x"21",x"AA",x"5C",x"0E",x"05",x"7E",x"8F",x"27",x"77",x"2B",x"0D",
x"20",x"F8",x"10",x"E7",x"AF",x"21",x"A6",x"5C",x"11",x"A1",x"5C",x"06",x"09",x"ED",x"6F",x"0E",
x"FF",x"ED",x"6F",x"20",x"04",x"0D",x"0C",x"20",x"0A",x"12",x"13",x"FD",x"34",x"71",x"FD",x"34",
x"72",x"0E",x"00",x"CB",x"40",x"28",x"01",x"23",x"10",x"E7",x"3A",x"AB",x"5C",x"D6",x"09",x"38",
x"0A",x"FD",x"35",x"71",x"3E",x"04",x"FD",x"BE",x"6F",x"18",x"41",x"EF",x"02",x"E2",x"38",x"EB",
x"CD",x"BA",x"2F",x"D9",x"3E",x"80",x"95",x"2E",x"00",x"CB",x"FA",x"D9",x"CD",x"DD",x"2F",x"FD",
x"7E",x"71",x"FE",x"08",x"38",x"06",x"D9",x"CB",x"12",x"D9",x"18",x"20",x"01",x"00",x"02",x"7B",
x"CD",x"8B",x"2F",x"5F",x"7A",x"CD",x"8B",x"2F",x"57",x"C5",x"D9",x"C1",x"10",x"F1",x"21",x"A1",
x"5C",x"79",x"FD",x"4E",x"71",x"09",x"77",x"FD",x"34",x"71",x"18",x"D3",x"F5",x"21",x"A1",x"5C",
x"FD",x"4E",x"71",x"06",x"00",x"09",x"41",x"F1",x"2B",x"7E",x"CE",x"00",x"77",x"A7",x"28",x"05",
x"FE",x"0A",x"3F",x"30",x"08",x"10",x"F1",x"36",x"01",x"04",x"FD",x"34",x"72",x"FD",x"70",x"71",
x"EF",x"02",x"38",x"D9",x"E1",x"D9",x"ED",x"4B",x"AB",x"5C",x"21",x"A1",x"5C",x"78",x"FE",x"09",
x"38",x"04",x"FE",x"FC",x"38",x"26",x"A7",x"CC",x"EF",x"15",x"AF",x"90",x"FA",x"52",x"2F",x"47",
x"18",x"0C",x"79",x"A7",x"28",x"03",x"7E",x"23",x"0D",x"CD",x"EF",x"15",x"10",x"F4",x"79",x"A7",
x"C8",x"04",x"3E",x"2E",x"D7",x"3E",x"30",x"10",x"FB",x"41",x"18",x"E6",x"50",x"15",x"06",x"01",
x"CD",x"4A",x"2F",x"3E",x"45",x"D7",x"4A",x"79",x"A7",x"F2",x"83",x"2F",x"ED",x"44",x"4F",x"3E",
x"2D",x"18",x"02",x"3E",x"2B",x"D7",x"06",x"00",x"C3",x"1B",x"1A",x"D5",x"6F",x"26",x"00",x"5D",
x"54",x"29",x"29",x"19",x"29",x"59",x"19",x"4C",x"7D",x"D1",x"C9",x"7E",x"36",x"00",x"A7",x"C8",
x"23",x"CB",x"7E",x"CB",x"FE",x"2B",x"C8",x"C5",x"01",x"05",x"00",x"09",x"41",x"4F",x"37",x"2B",
x"7E",x"2F",x"CE",x"00",x"77",x"10",x"F8",x"79",x"C1",x"C9",x"E5",x"F5",x"4E",x"23",x"46",x"77",
x"23",x"79",x"4E",x"C5",x"23",x"4E",x"23",x"46",x"EB",x"57",x"5E",x"D5",x"23",x"56",x"23",x"5E",
x"D5",x"D9",x"D1",x"E1",x"C1",x"D9",x"23",x"56",x"23",x"5E",x"F1",x"E1",x"C9",x"A7",x"C8",x"FE",
x"21",x"30",x"16",x"C5",x"47",x"D9",x"CB",x"2D",x"CB",x"1A",x"CB",x"1B",x"D9",x"CB",x"1A",x"CB",
x"1B",x"10",x"F2",x"C1",x"D0",x"CD",x"04",x"30",x"C0",x"D9",x"AF",x"2E",x"00",x"57",x"5D",x"D9",
x"11",x"00",x"00",x"C9",x"1C",x"C0",x"14",x"C0",x"D9",x"1C",x"20",x"01",x"14",x"D9",x"C9",x"EB",
x"CD",x"6E",x"34",x"EB",x"1A",x"B6",x"20",x"26",x"D5",x"23",x"E5",x"23",x"5E",x"23",x"56",x"23",
x"23",x"23",x"7E",x"23",x"4E",x"23",x"46",x"E1",x"EB",x"09",x"EB",x"8E",x"0F",x"CE",x"00",x"20",
x"0B",x"9F",x"77",x"23",x"73",x"23",x"72",x"2B",x"2B",x"2B",x"D1",x"C9",x"2B",x"D1",x"CD",x"93",
x"32",x"D9",x"E5",x"D9",x"D5",x"E5",x"CD",x"9B",x"2F",x"47",x"EB",x"CD",x"9B",x"2F",x"4F",x"B8",
x"30",x"03",x"78",x"41",x"EB",x"F5",x"90",x"CD",x"BA",x"2F",x"CD",x"DD",x"2F",x"F1",x"E1",x"77",
x"E5",x"68",x"61",x"19",x"D9",x"EB",x"ED",x"4A",x"EB",x"7C",x"8D",x"6F",x"1F",x"AD",x"D9",x"EB",
x"E1",x"1F",x"30",x"08",x"3E",x"01",x"CD",x"DD",x"2F",x"34",x"28",x"23",x"D9",x"7D",x"E6",x"80",
x"D9",x"23",x"77",x"2B",x"28",x"1F",x"7B",x"ED",x"44",x"3F",x"5F",x"7A",x"2F",x"CE",x"00",x"57",
x"D9",x"7B",x"2F",x"CE",x"00",x"5F",x"7A",x"2F",x"CE",x"00",x"30",x"07",x"1F",x"D9",x"34",x"CA",
x"AD",x"31",x"D9",x"57",x"D9",x"AF",x"C3",x"55",x"31",x"C5",x"06",x"10",x"7C",x"4D",x"21",x"00",
x"00",x"29",x"38",x"0A",x"CB",x"11",x"17",x"30",x"03",x"19",x"38",x"02",x"10",x"F3",x"C1",x"C9",
x"CD",x"E9",x"34",x"D8",x"23",x"AE",x"CB",x"FE",x"2B",x"C9",x"1A",x"B6",x"20",x"22",x"D5",x"E5",
x"D5",x"CD",x"7F",x"2D",x"EB",x"E3",x"41",x"CD",x"7F",x"2D",x"78",x"A9",x"4F",x"E1",x"CD",x"A9",
x"30",x"EB",x"E1",x"38",x"0A",x"7A",x"B3",x"20",x"01",x"4F",x"CD",x"8E",x"2D",x"D1",x"C9",x"D1",
x"CD",x"93",x"32",x"AF",x"CD",x"C0",x"30",x"D8",x"D9",x"E5",x"D9",x"D5",x"EB",x"CD",x"C0",x"30",
x"EB",x"38",x"5A",x"E5",x"CD",x"BA",x"2F",x"78",x"A7",x"ED",x"62",x"D9",x"E5",x"ED",x"62",x"D9",
x"06",x"21",x"18",x"11",x"30",x"05",x"19",x"D9",x"ED",x"5A",x"D9",x"D9",x"CB",x"1C",x"CB",x"1D",
x"D9",x"CB",x"1C",x"CB",x"1D",x"D9",x"CB",x"18",x"CB",x"19",x"D9",x"CB",x"19",x"1F",x"10",x"E4",
x"EB",x"D9",x"EB",x"D9",x"C1",x"E1",x"78",x"81",x"20",x"01",x"A7",x"3D",x"3F",x"17",x"3F",x"1F",
x"F2",x"46",x"31",x"30",x"68",x"A7",x"3C",x"20",x"08",x"38",x"06",x"D9",x"CB",x"7A",x"D9",x"20",
x"5C",x"77",x"D9",x"78",x"D9",x"30",x"15",x"7E",x"A7",x"3E",x"80",x"28",x"01",x"AF",x"D9",x"A2",
x"CD",x"FB",x"2F",x"07",x"77",x"38",x"2E",x"23",x"77",x"2B",x"18",x"29",x"06",x"20",x"D9",x"CB",
x"7A",x"D9",x"20",x"12",x"07",x"CB",x"13",x"CB",x"12",x"D9",x"CB",x"13",x"CB",x"12",x"D9",x"35",
x"28",x"D7",x"10",x"EA",x"18",x"D7",x"17",x"30",x"0C",x"CD",x"04",x"30",x"20",x"07",x"D9",x"16",
x"80",x"D9",x"34",x"28",x"18",x"E5",x"23",x"D9",x"D5",x"D9",x"C1",x"78",x"17",x"CB",x"16",x"1F",
x"77",x"23",x"71",x"23",x"72",x"23",x"73",x"E1",x"D1",x"D9",x"E1",x"D9",x"C9",x"CF",x"05",x"CD",
x"93",x"32",x"EB",x"AF",x"CD",x"C0",x"30",x"38",x"F4",x"EB",x"CD",x"C0",x"30",x"D8",x"D9",x"E5",
x"D9",x"D5",x"E5",x"CD",x"BA",x"2F",x"D9",x"E5",x"60",x"69",x"D9",x"61",x"68",x"AF",x"06",x"DF",
x"18",x"10",x"17",x"CB",x"11",x"D9",x"CB",x"11",x"CB",x"10",x"D9",x"29",x"D9",x"ED",x"6A",x"D9",
x"38",x"10",x"ED",x"52",x"D9",x"ED",x"52",x"D9",x"30",x"0F",x"19",x"D9",x"ED",x"5A",x"D9",x"A7",
x"18",x"08",x"A7",x"ED",x"52",x"D9",x"ED",x"52",x"D9",x"37",x"04",x"FA",x"D2",x"31",x"F5",x"28",
x"E1",x"5F",x"51",x"D9",x"59",x"50",x"F1",x"CB",x"18",x"F1",x"CB",x"18",x"D9",x"C1",x"E1",x"78",
x"91",x"C3",x"3D",x"31",x"7E",x"A7",x"C8",x"FE",x"81",x"30",x"06",x"36",x"00",x"3E",x"20",x"18",
x"51",x"FE",x"91",x"20",x"1A",x"23",x"23",x"23",x"3E",x"80",x"A6",x"2B",x"B6",x"2B",x"20",x"03",
x"3E",x"80",x"AE",x"2B",x"20",x"36",x"77",x"23",x"36",x"FF",x"2B",x"3E",x"18",x"18",x"33",x"30",
x"2C",x"D5",x"2F",x"C6",x"91",x"23",x"56",x"23",x"5E",x"2B",x"2B",x"0E",x"00",x"CB",x"7A",x"28",
x"01",x"0D",x"CB",x"FA",x"06",x"08",x"90",x"80",x"38",x"04",x"5A",x"16",x"00",x"90",x"28",x"07",
x"47",x"CB",x"3A",x"CB",x"1B",x"10",x"FA",x"CD",x"8E",x"2D",x"D1",x"C9",x"7E",x"D6",x"A0",x"F0",
x"ED",x"44",x"D5",x"EB",x"2B",x"47",x"CB",x"38",x"CB",x"38",x"CB",x"38",x"28",x"05",x"36",x"00",
x"2B",x"10",x"FB",x"E6",x"07",x"28",x"09",x"47",x"3E",x"FF",x"CB",x"27",x"10",x"FC",x"A6",x"77",
x"EB",x"D1",x"C9",x"CD",x"96",x"32",x"EB",x"7E",x"A7",x"C0",x"D5",x"CD",x"7F",x"2D",x"AF",x"23",
x"77",x"2B",x"77",x"06",x"91",x"7A",x"A7",x"20",x"08",x"B3",x"42",x"28",x"10",x"53",x"58",x"06",
x"89",x"EB",x"05",x"29",x"30",x"FC",x"CB",x"09",x"CB",x"1C",x"CB",x"1D",x"EB",x"2B",x"73",x"2B",
x"72",x"2B",x"70",x"D1",x"C9",x"00",x"B0",x"00",x"40",x"B0",x"00",x"01",x"30",x"00",x"F1",x"49",
x"0F",x"DA",x"A2",x"40",x"B0",x"00",x"0A",x"8F",x"36",x"3C",x"34",x"A1",x"33",x"0F",x"30",x"CA",
x"30",x"AF",x"31",x"51",x"38",x"1B",x"35",x"24",x"35",x"3B",x"35",x"3B",x"35",x"3B",x"35",x"3B",
x"35",x"3B",x"35",x"3B",x"35",x"14",x"30",x"2D",x"35",x"3B",x"35",x"3B",x"35",x"3B",x"35",x"3B",
x"35",x"3B",x"35",x"3B",x"35",x"9C",x"35",x"DE",x"35",x"BC",x"34",x"45",x"36",x"6E",x"34",x"69",
x"36",x"DE",x"35",x"74",x"36",x"B5",x"37",x"AA",x"37",x"DA",x"37",x"33",x"38",x"43",x"38",x"E2",
x"37",x"13",x"37",x"C4",x"36",x"AF",x"36",x"4A",x"38",x"92",x"34",x"6A",x"34",x"AC",x"34",x"A5",
x"34",x"B3",x"34",x"1F",x"36",x"C9",x"35",x"01",x"35",x"C0",x"33",x"A0",x"36",x"86",x"36",x"C6",
x"33",x"7A",x"36",x"06",x"35",x"F9",x"34",x"9B",x"36",x"83",x"37",x"14",x"32",x"A2",x"33",x"4F",
x"2D",x"97",x"32",x"49",x"34",x"1B",x"34",x"2D",x"34",x"0F",x"34",x"CD",x"BF",x"35",x"78",x"32",
x"67",x"5C",x"D9",x"E3",x"D9",x"ED",x"53",x"65",x"5C",x"D9",x"7E",x"23",x"E5",x"A7",x"F2",x"80",
x"33",x"57",x"E6",x"60",x"0F",x"0F",x"0F",x"0F",x"C6",x"7C",x"6F",x"7A",x"E6",x"1F",x"18",x"0E",
x"FE",x"18",x"30",x"08",x"D9",x"01",x"FB",x"FF",x"54",x"5D",x"09",x"D9",x"07",x"6F",x"11",x"D7",
x"32",x"26",x"00",x"19",x"5E",x"23",x"56",x"21",x"65",x"33",x"E3",x"D5",x"D9",x"ED",x"4B",x"66",
x"5C",x"C9",x"F1",x"3A",x"67",x"5C",x"D9",x"18",x"C3",x"D5",x"E5",x"01",x"05",x"00",x"CD",x"05",
x"1F",x"E1",x"D1",x"C9",x"ED",x"5B",x"65",x"5C",x"CD",x"C0",x"33",x"ED",x"53",x"65",x"5C",x"C9",
x"CD",x"A9",x"33",x"ED",x"B0",x"C9",x"62",x"6B",x"CD",x"A9",x"33",x"D9",x"E5",x"D9",x"E3",x"C5",
x"7E",x"E6",x"C0",x"07",x"07",x"4F",x"0C",x"7E",x"E6",x"3F",x"20",x"02",x"23",x"7E",x"C6",x"50",
x"12",x"3E",x"05",x"91",x"23",x"13",x"06",x"00",x"ED",x"B0",x"C1",x"E3",x"D9",x"E1",x"D9",x"47",
x"AF",x"05",x"C8",x"12",x"13",x"18",x"FA",x"A7",x"C8",x"F5",x"D5",x"11",x"00",x"00",x"CD",x"C8",
x"33",x"D1",x"F1",x"3D",x"18",x"F2",x"4F",x"07",x"07",x"81",x"4F",x"06",x"00",x"09",x"C9",x"D5",
x"2A",x"68",x"5C",x"CD",x"06",x"34",x"CD",x"C0",x"33",x"E1",x"C9",x"62",x"6B",x"D9",x"E5",x"21",
x"C5",x"32",x"D9",x"CD",x"F7",x"33",x"CD",x"C8",x"33",x"D9",x"E1",x"D9",x"C9",x"E5",x"EB",x"2A",
x"68",x"5C",x"CD",x"06",x"34",x"EB",x"CD",x"C0",x"33",x"EB",x"E1",x"C9",x"06",x"05",x"1A",x"4E",
x"EB",x"12",x"71",x"23",x"13",x"10",x"F7",x"EB",x"C9",x"47",x"CD",x"5E",x"33",x"31",x"0F",x"C0",
x"02",x"A0",x"C2",x"31",x"E0",x"04",x"E2",x"C1",x"03",x"38",x"CD",x"C6",x"33",x"CD",x"62",x"33",
x"0F",x"01",x"C2",x"02",x"35",x"EE",x"E1",x"03",x"38",x"C9",x"06",x"FF",x"18",x"06",x"CD",x"E9",
x"34",x"D8",x"06",x"00",x"7E",x"A7",x"28",x"0B",x"23",x"78",x"E6",x"80",x"B6",x"17",x"3F",x"1F",
x"77",x"2B",x"C9",x"D5",x"E5",x"CD",x"7F",x"2D",x"E1",x"78",x"B1",x"2F",x"4F",x"CD",x"8E",x"2D",
x"D1",x"C9",x"CD",x"E9",x"34",x"D8",x"D5",x"11",x"01",x"00",x"23",x"CB",x"16",x"2B",x"9F",x"4F",
x"CD",x"8E",x"2D",x"D1",x"C9",x"CD",x"99",x"1E",x"ED",x"78",x"18",x"04",x"CD",x"99",x"1E",x"0A",
x"C3",x"28",x"2D",x"CD",x"99",x"1E",x"21",x"2B",x"2D",x"E5",x"C5",x"C9",x"CD",x"F1",x"2B",x"0B",
x"78",x"B1",x"20",x"23",x"1A",x"CD",x"8D",x"2C",x"38",x"09",x"D6",x"90",x"38",x"19",x"FE",x"15",
x"30",x"15",x"3C",x"3D",x"87",x"87",x"87",x"FE",x"A8",x"30",x"0C",x"ED",x"4B",x"7B",x"5C",x"81",
x"4F",x"30",x"01",x"04",x"C3",x"2B",x"2D",x"CF",x"09",x"E5",x"C5",x"47",x"7E",x"23",x"B6",x"23",
x"B6",x"23",x"B6",x"78",x"C1",x"E1",x"C0",x"37",x"C9",x"CD",x"E9",x"34",x"D8",x"3E",x"FF",x"18",
x"06",x"CD",x"E9",x"34",x"18",x"05",x"AF",x"23",x"AE",x"2B",x"07",x"E5",x"3E",x"00",x"77",x"23",
x"77",x"23",x"17",x"77",x"1F",x"23",x"77",x"23",x"77",x"E1",x"C9",x"EB",x"CD",x"E9",x"34",x"EB",
x"D8",x"37",x"18",x"E7",x"EB",x"CD",x"E9",x"34",x"EB",x"D0",x"A7",x"18",x"DE",x"EB",x"CD",x"E9",
x"34",x"EB",x"D0",x"D5",x"1B",x"AF",x"12",x"1B",x"12",x"D1",x"C9",x"78",x"D6",x"08",x"CB",x"57",
x"20",x"01",x"3D",x"0F",x"30",x"08",x"F5",x"E5",x"CD",x"3C",x"34",x"D1",x"EB",x"F1",x"CB",x"57",
x"20",x"07",x"0F",x"F5",x"CD",x"0F",x"30",x"18",x"33",x"0F",x"F5",x"CD",x"F1",x"2B",x"D5",x"C5",
x"CD",x"F1",x"2B",x"E1",x"7C",x"B5",x"E3",x"78",x"20",x"0B",x"B1",x"C1",x"28",x"04",x"F1",x"3F",
x"18",x"16",x"F1",x"18",x"13",x"B1",x"28",x"0D",x"1A",x"96",x"38",x"09",x"20",x"ED",x"0B",x"13",
x"23",x"E3",x"2B",x"18",x"DF",x"C1",x"F1",x"A7",x"F5",x"EF",x"A0",x"38",x"F1",x"F5",x"DC",x"01",
x"35",x"F1",x"F5",x"D4",x"F9",x"34",x"F1",x"0F",x"D4",x"01",x"35",x"C9",x"CD",x"F1",x"2B",x"D5",
x"C5",x"CD",x"F1",x"2B",x"E1",x"E5",x"D5",x"C5",x"09",x"44",x"4D",x"F7",x"CD",x"B2",x"2A",x"C1",
x"E1",x"78",x"B1",x"28",x"02",x"ED",x"B0",x"C1",x"E1",x"78",x"B1",x"28",x"02",x"ED",x"B0",x"2A",
x"65",x"5C",x"11",x"FB",x"FF",x"E5",x"19",x"D1",x"C9",x"CD",x"D5",x"2D",x"38",x"0E",x"20",x"0C",
x"F5",x"01",x"01",x"00",x"F7",x"F1",x"12",x"CD",x"B2",x"2A",x"EB",x"C9",x"CF",x"0A",x"2A",x"5D",
x"5C",x"E5",x"78",x"C6",x"E3",x"9F",x"F5",x"CD",x"F1",x"2B",x"D5",x"03",x"F7",x"E1",x"ED",x"53",
x"5D",x"5C",x"D5",x"ED",x"B0",x"EB",x"2B",x"36",x"0D",x"FD",x"CB",x"01",x"BE",x"CD",x"FB",x"24",
x"DF",x"FE",x"0D",x"20",x"07",x"E1",x"F1",x"FD",x"AE",x"01",x"E6",x"40",x"C2",x"8A",x"1C",x"22",
x"5D",x"5C",x"FD",x"CB",x"01",x"FE",x"CD",x"FB",x"24",x"E1",x"22",x"5D",x"5C",x"18",x"A0",x"01",
x"01",x"00",x"F7",x"22",x"5B",x"5C",x"E5",x"2A",x"51",x"5C",x"E5",x"3E",x"FF",x"CD",x"01",x"16",
x"CD",x"E3",x"2D",x"E1",x"CD",x"15",x"16",x"D1",x"2A",x"5B",x"5C",x"A7",x"ED",x"52",x"44",x"4D",
x"CD",x"B2",x"2A",x"EB",x"C9",x"CD",x"94",x"1E",x"FE",x"10",x"D2",x"9F",x"1E",x"2A",x"51",x"5C",
x"E5",x"CD",x"01",x"16",x"CD",x"E6",x"15",x"01",x"00",x"00",x"30",x"03",x"0C",x"F7",x"12",x"CD",
x"B2",x"2A",x"E1",x"CD",x"15",x"16",x"C3",x"BF",x"35",x"CD",x"F1",x"2B",x"78",x"B1",x"28",x"01",
x"1A",x"C3",x"28",x"2D",x"CD",x"F1",x"2B",x"C3",x"2B",x"2D",x"D9",x"E5",x"21",x"67",x"5C",x"35",
x"E1",x"20",x"04",x"23",x"D9",x"C9",x"D9",x"5E",x"7B",x"17",x"9F",x"57",x"19",x"D9",x"C9",x"13",
x"13",x"1A",x"1B",x"1B",x"A7",x"20",x"EF",x"D9",x"23",x"D9",x"C9",x"F1",x"D9",x"E3",x"D9",x"C9",
x"EF",x"C0",x"02",x"31",x"E0",x"05",x"27",x"E0",x"01",x"C0",x"04",x"03",x"E0",x"38",x"C9",x"EF",
x"31",x"36",x"00",x"04",x"3A",x"38",x"C9",x"31",x"3A",x"C0",x"03",x"E0",x"01",x"30",x"00",x"03",
x"A1",x"03",x"38",x"C9",x"EF",x"3D",x"34",x"F1",x"38",x"AA",x"3B",x"29",x"04",x"31",x"27",x"C3",
x"03",x"31",x"0F",x"A1",x"03",x"88",x"13",x"36",x"58",x"65",x"66",x"9D",x"78",x"65",x"40",x"A2",
x"60",x"32",x"C9",x"E7",x"21",x"F7",x"AF",x"24",x"EB",x"2F",x"B0",x"B0",x"14",x"EE",x"7E",x"BB",
x"94",x"58",x"F1",x"3A",x"7E",x"F8",x"CF",x"E3",x"38",x"CD",x"D5",x"2D",x"20",x"07",x"38",x"03",
x"86",x"30",x"09",x"CF",x"05",x"38",x"07",x"96",x"30",x"04",x"ED",x"44",x"77",x"C9",x"EF",x"02",
x"A0",x"38",x"C9",x"EF",x"3D",x"31",x"37",x"00",x"04",x"38",x"CF",x"09",x"A0",x"02",x"38",x"7E",
x"36",x"80",x"CD",x"28",x"2D",x"EF",x"34",x"38",x"00",x"03",x"01",x"31",x"34",x"F0",x"4C",x"CC",
x"CC",x"CD",x"03",x"37",x"00",x"08",x"01",x"A1",x"03",x"01",x"38",x"34",x"EF",x"01",x"34",x"F0",
x"31",x"72",x"17",x"F8",x"04",x"01",x"A2",x"03",x"A2",x"03",x"31",x"34",x"32",x"20",x"04",x"A2",
x"03",x"8C",x"11",x"AC",x"14",x"09",x"56",x"DA",x"A5",x"59",x"30",x"C5",x"5C",x"90",x"AA",x"9E",
x"70",x"6F",x"61",x"A1",x"CB",x"DA",x"96",x"A4",x"31",x"9F",x"B4",x"E7",x"A0",x"FE",x"5C",x"FC",
x"EA",x"1B",x"43",x"CA",x"36",x"ED",x"A7",x"9C",x"7E",x"5E",x"F0",x"6E",x"23",x"80",x"93",x"04",
x"0F",x"38",x"C9",x"EF",x"3D",x"34",x"EE",x"22",x"F9",x"83",x"6E",x"04",x"31",x"A2",x"0F",x"27",
x"03",x"31",x"0F",x"31",x"0F",x"31",x"2A",x"A1",x"03",x"31",x"37",x"C0",x"00",x"04",x"02",x"38",
x"C9",x"A1",x"03",x"01",x"36",x"00",x"02",x"1B",x"38",x"C9",x"EF",x"39",x"2A",x"A1",x"03",x"E0",
x"00",x"06",x"1B",x"33",x"03",x"EF",x"39",x"31",x"31",x"04",x"31",x"0F",x"A1",x"03",x"86",x"14",
x"E6",x"5C",x"1F",x"0B",x"A3",x"8F",x"38",x"EE",x"E9",x"15",x"63",x"BB",x"23",x"EE",x"92",x"0D",
x"CD",x"ED",x"F1",x"23",x"5D",x"1B",x"EA",x"04",x"38",x"C9",x"EF",x"31",x"1F",x"01",x"20",x"05",
x"38",x"C9",x"CD",x"97",x"32",x"7E",x"FE",x"81",x"38",x"0E",x"EF",x"A1",x"1B",x"01",x"05",x"31",
x"36",x"A3",x"01",x"00",x"06",x"1B",x"33",x"03",x"EF",x"A0",x"01",x"31",x"31",x"04",x"31",x"0F",
x"A1",x"03",x"8C",x"10",x"B2",x"13",x"0E",x"55",x"E4",x"8D",x"58",x"39",x"BC",x"5B",x"98",x"FD",
x"9E",x"00",x"36",x"75",x"A0",x"DB",x"E8",x"B4",x"63",x"42",x"C4",x"E6",x"B5",x"09",x"36",x"BE",
x"E9",x"36",x"73",x"1B",x"5D",x"EC",x"D8",x"DE",x"63",x"BE",x"F0",x"61",x"A1",x"B3",x"0C",x"04",
x"0F",x"38",x"C9",x"EF",x"31",x"31",x"04",x"A1",x"03",x"1B",x"28",x"A1",x"0F",x"05",x"24",x"31",
x"0F",x"38",x"C9",x"EF",x"22",x"A3",x"03",x"1B",x"38",x"C9",x"EF",x"31",x"30",x"00",x"1E",x"A2",
x"38",x"EF",x"01",x"31",x"30",x"00",x"07",x"25",x"04",x"38",x"C3",x"C4",x"36",x"02",x"31",x"30",
x"00",x"09",x"A0",x"01",x"37",x"00",x"06",x"A1",x"01",x"05",x"02",x"A1",x"38",x"C9",x"FF",x"FF",
x"F6",x"20",x"FE",x"6E",x"C2",x"C4",x"0C",x"21",x"BF",x"04",x"CB",x"46",x"28",x"0D",x"CB",x"86",
x"3E",x"04",x"CD",x"B7",x"0E",x"CD",x"B5",x"0E",x"CD",x"B5",x"0E",x"C3",x"00",x"0D",x"C3",x"CB",
x"11",x"3E",x"02",x"CD",x"01",x"16",x"2A",x"5D",x"5C",x"CD",x"71",x"3B",x"FE",x"0D",x"CA",x"B2",
x"1B",x"11",x"7A",x"3B",x"CD",x"60",x"3B",x"CA",x"A4",x"3A",x"11",x"7E",x"3B",x"CD",x"60",x"3B",
x"CA",x"E3",x"39",x"11",x"83",x"3B",x"CD",x"60",x"3B",x"CA",x"32",x"3A",x"3E",x"15",x"CD",x"B7",
x"0E",x"7E",x"23",x"FE",x"0D",x"28",x"03",x"B7",x"20",x"F4",x"AF",x"CD",x"B7",x"0E",x"CD",x"B5",
x"0E",x"FE",x"02",x"28",x"13",x"FE",x"05",x"28",x"15",x"FE",x"09",x"28",x"19",x"FE",x"0A",x"28",
x"24",x"FE",x"0B",x"28",x"0C",x"C3",x"1D",x"39",x"CD",x"2D",x"39",x"CD",x"B5",x"0E",x"C3",x"B2",
x"1B",x"CD",x"2D",x"39",x"18",x"D8",x"CD",x"14",x"39",x"7E",x"CD",x"B7",x"0E",x"23",x"1B",x"7A",
x"B3",x"20",x"F6",x"18",x"C9",x"CD",x"14",x"39",x"CD",x"B5",x"0E",x"77",x"23",x"1B",x"7A",x"B3",
x"20",x"F6",x"18",x"BA",x"CD",x"AD",x"39",x"EB",x"CD",x"AD",x"39",x"EB",x"C9",x"3E",x"02",x"D3",
x"FE",x"21",x"88",x"3B",x"7E",x"B7",x"CA",x"B2",x"1B",x"D7",x"23",x"18",x"F7",x"21",x"BF",x"04",
x"36",x"01",x"CD",x"B5",x"0E",x"B7",x"28",x"03",x"D7",x"18",x"F7",x"21",x"BF",x"04",x"36",x"00",
x"C9",x"09",x"CD",x"71",x"3B",x"B7",x"C8",x"FE",x"0D",x"C9",x"3E",x"11",x"CD",x"B7",x"0E",x"7E",
x"FE",x"0D",x"28",x"06",x"B7",x"28",x"03",x"23",x"18",x"F2",x"AF",x"CD",x"B7",x"0E",x"CD",x"B5",
x"0E",x"FE",x"7F",x"28",x"2A",x"FE",x"80",x"C9",x"3E",x"10",x"CD",x"B7",x"0E",x"7E",x"FE",x"0D",
x"28",x"06",x"B7",x"28",x"03",x"23",x"18",x"F2",x"AF",x"CD",x"B7",x"0E",x"CD",x"B5",x"0E",x"FE",
x"7F",x"28",x"0C",x"CD",x"AD",x"39",x"22",x"B8",x"04",x"CD",x"B5",x"0E",x"FE",x"80",x"C9",x"3E",
x"01",x"B7",x"C9",x"3E",x"13",x"CD",x"B7",x"0E",x"AF",x"CD",x"B7",x"0E",x"3E",x"02",x"CD",x"B7",
x"0E",x"CD",x"B5",x"0E",x"4F",x"CD",x"B5",x"0E",x"47",x"CD",x"B5",x"0E",x"C9",x"CD",x"B5",x"0E",
x"6F",x"CD",x"B5",x"0E",x"67",x"C9",x"2A",x"59",x"5C",x"ED",x"5B",x"53",x"5C",x"37",x"ED",x"52",
x"44",x"4D",x"2A",x"4B",x"5C",x"ED",x"52",x"EB",x"C9",x"3E",x"14",x"CD",x"B7",x"0E",x"AF",x"CD",
x"B7",x"0E",x"3E",x"02",x"CD",x"B7",x"0E",x"79",x"CD",x"B7",x"0E",x"78",x"CD",x"B7",x"0E",x"CD",
x"B5",x"0E",x"C9",x"01",x"04",x"00",x"CD",x"41",x"39",x"CA",x"1D",x"39",x"CD",x"4A",x"39",x"C2",
x"1D",x"39",x"CD",x"B6",x"39",x"C5",x"CD",x"C9",x"39",x"42",x"4B",x"CD",x"C9",x"39",x"C1",x"3E",
x"14",x"CD",x"B7",x"0E",x"79",x"CD",x"B7",x"0E",x"78",x"CD",x"B7",x"0E",x"7E",x"CD",x"B7",x"0E",
x"23",x"0B",x"78",x"B1",x"20",x"F6",x"CD",x"B5",x"0E",x"3E",x"12",x"CD",x"B7",x"0E",x"CD",x"B5",
x"0E",x"C3",x"B2",x"1B",x"3E",x"13",x"CD",x"B7",x"0E",x"7B",x"CD",x"B7",x"0E",x"7A",x"CD",x"B7",
x"0E",x"C9",x"01",x"04",x"00",x"CD",x"41",x"39",x"CA",x"1D",x"39",x"CD",x"68",x"39",x"C2",x"1D",
x"39",x"CD",x"93",x"39",x"ED",x"43",x"B0",x"04",x"CD",x"93",x"39",x"ED",x"43",x"B2",x"04",x"CD",
x"B6",x"39",x"50",x"59",x"2A",x"B0",x"04",x"37",x"ED",x"52",x"38",x"09",x"11",x"05",x"00",x"19",
x"44",x"4D",x"CD",x"05",x"1F",x"CD",x"B6",x"39",x"EB",x"2A",x"59",x"5C",x"2B",x"ED",x"4B",x"B0",
x"04",x"C5",x"CD",x"E5",x"19",x"C1",x"E5",x"C5",x"CD",x"55",x"16",x"23",x"ED",x"4B",x"B2",x"04",
x"09",x"22",x"4B",x"5C",x"D1",x"E1",x"CD",x"24",x"3A",x"CD",x"B5",x"0E",x"77",x"23",x"1B",x"7A",
x"B3",x"20",x"F6",x"CD",x"B5",x"0E",x"C3",x"19",x"3A",x"3E",x"12",x"CD",x"B7",x"0E",x"CD",x"B5",
x"0E",x"C3",x"1D",x"39",x"01",x"03",x"00",x"CD",x"41",x"39",x"CA",x"1D",x"39",x"CD",x"68",x"39",
x"C2",x"1D",x"39",x"2A",x"B8",x"04",x"11",x"1B",x"C0",x"B7",x"ED",x"52",x"C2",x"1D",x"39",x"CD",
x"24",x"3A",x"F3",x"CD",x"B5",x"0E",x"ED",x"47",x"CD",x"AD",x"39",x"E5",x"CD",x"AD",x"39",x"EB",
x"CD",x"AD",x"39",x"44",x"4D",x"CD",x"AD",x"39",x"E5",x"F1",x"08",x"E1",x"D9",x"CD",x"AD",x"39",
x"22",x"B4",x"04",x"CD",x"AD",x"39",x"EB",x"CD",x"AD",x"39",x"44",x"4D",x"CD",x"AD",x"39",x"E5",
x"FD",x"E1",x"CD",x"AD",x"39",x"E5",x"DD",x"E1",x"CD",x"B5",x"0E",x"E6",x"02",x"0F",x"32",x"B0",
x"04",x"CD",x"B5",x"0E",x"ED",x"4F",x"31",x"BE",x"04",x"CD",x"AD",x"39",x"E5",x"CD",x"AD",x"39",
x"22",x"B2",x"04",x"CD",x"B5",x"0E",x"A7",x"28",x"07",x"3D",x"28",x"08",x"ED",x"5E",x"18",x"06",
x"ED",x"46",x"18",x"02",x"ED",x"56",x"CD",x"B5",x"0E",x"E6",x"07",x"F5",x"21",x"00",x"40",x"CD",
x"B5",x"0E",x"77",x"E6",x"07",x"D3",x"FE",x"23",x"7C",x"B5",x"20",x"F3",x"CD",x"B5",x"0E",x"3E",
x"12",x"CD",x"B7",x"0E",x"CD",x"B5",x"0E",x"F1",x"D3",x"FE",x"2A",x"B4",x"04",x"3A",x"B0",x"04",
x"0F",x"38",x"06",x"F1",x"ED",x"7B",x"B2",x"04",x"C9",x"F1",x"ED",x"7B",x"B2",x"04",x"FB",x"C9",
x"E5",x"D5",x"1A",x"FE",x"00",x"28",x"07",x"BE",x"20",x"04",x"23",x"13",x"18",x"F4",x"D1",x"E1",
x"C9",x"3E",x"20",x"2B",x"23",x"BE",x"28",x"FC",x"7E",x"C9",x"73",x"6E",x"61",x"00",x"73",x"61",
x"76",x"65",x"00",x"6C",x"6F",x"61",x"64",x"00",x"49",x"2F",x"4F",x"20",x"45",x"72",x"72",x"6F",
x"72",x"2E",x"0D",x"00",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",x"FF",
x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"10",x"10",x"10",x"10",x"00",x"10",x"00",
x"00",x"24",x"24",x"00",x"00",x"00",x"00",x"00",x"00",x"24",x"7E",x"24",x"24",x"7E",x"24",x"00",
x"00",x"08",x"3E",x"28",x"3E",x"0A",x"3E",x"08",x"00",x"62",x"64",x"08",x"10",x"26",x"46",x"00",
x"00",x"10",x"28",x"10",x"2A",x"44",x"3A",x"00",x"00",x"08",x"10",x"00",x"00",x"00",x"00",x"00",
x"00",x"04",x"08",x"08",x"08",x"08",x"04",x"00",x"00",x"20",x"10",x"10",x"10",x"10",x"20",x"00",
x"00",x"00",x"14",x"08",x"3E",x"08",x"14",x"00",x"00",x"00",x"08",x"08",x"3E",x"08",x"08",x"00",
x"00",x"00",x"00",x"00",x"00",x"08",x"08",x"10",x"00",x"00",x"00",x"00",x"3E",x"00",x"00",x"00",
x"00",x"00",x"00",x"00",x"00",x"18",x"18",x"00",x"00",x"00",x"02",x"04",x"08",x"10",x"20",x"00",
x"00",x"3C",x"46",x"4A",x"52",x"62",x"3C",x"00",x"00",x"18",x"28",x"08",x"08",x"08",x"3E",x"00",
x"00",x"3C",x"42",x"02",x"3C",x"40",x"7E",x"00",x"00",x"3C",x"42",x"0C",x"02",x"42",x"3C",x"00",
x"00",x"08",x"18",x"28",x"48",x"7E",x"08",x"00",x"00",x"7E",x"40",x"7C",x"02",x"42",x"3C",x"00",
x"00",x"3C",x"40",x"7C",x"42",x"42",x"3C",x"00",x"00",x"7E",x"02",x"04",x"08",x"10",x"10",x"00",
x"00",x"3C",x"42",x"3C",x"42",x"42",x"3C",x"00",x"00",x"3C",x"42",x"42",x"3E",x"02",x"3C",x"00",
x"00",x"00",x"00",x"10",x"00",x"00",x"10",x"00",x"00",x"00",x"10",x"00",x"00",x"10",x"10",x"20",
x"00",x"00",x"04",x"08",x"10",x"08",x"04",x"00",x"00",x"00",x"00",x"3E",x"00",x"3E",x"00",x"00",
x"00",x"00",x"10",x"08",x"04",x"08",x"10",x"00",x"00",x"3C",x"42",x"04",x"08",x"00",x"08",x"00",
x"00",x"3C",x"4A",x"56",x"5E",x"40",x"3C",x"00",x"00",x"3C",x"42",x"42",x"7E",x"42",x"42",x"00",
x"00",x"7C",x"42",x"7C",x"42",x"42",x"7C",x"00",x"00",x"3C",x"42",x"40",x"40",x"42",x"3C",x"00",
x"00",x"78",x"44",x"42",x"42",x"44",x"78",x"00",x"00",x"7E",x"40",x"7C",x"40",x"40",x"7E",x"00",
x"00",x"7E",x"40",x"7C",x"40",x"40",x"40",x"00",x"00",x"3C",x"42",x"40",x"4E",x"42",x"3C",x"00",
x"00",x"42",x"42",x"7E",x"42",x"42",x"42",x"00",x"00",x"3E",x"08",x"08",x"08",x"08",x"3E",x"00",
x"00",x"02",x"02",x"02",x"42",x"42",x"3C",x"00",x"00",x"44",x"48",x"70",x"48",x"44",x"42",x"00",
x"00",x"40",x"40",x"40",x"40",x"40",x"7E",x"00",x"00",x"42",x"66",x"5A",x"42",x"42",x"42",x"00",
x"00",x"42",x"62",x"52",x"4A",x"46",x"42",x"00",x"00",x"3C",x"42",x"42",x"42",x"42",x"3C",x"00",
x"00",x"7C",x"42",x"42",x"7C",x"40",x"40",x"00",x"00",x"3C",x"42",x"42",x"52",x"4A",x"3C",x"00",
x"00",x"7C",x"42",x"42",x"7C",x"44",x"42",x"00",x"00",x"3C",x"40",x"3C",x"02",x"42",x"3C",x"00",
x"00",x"FE",x"10",x"10",x"10",x"10",x"10",x"00",x"00",x"42",x"42",x"42",x"42",x"42",x"3C",x"00",
x"00",x"42",x"42",x"42",x"42",x"24",x"18",x"00",x"00",x"42",x"42",x"42",x"42",x"5A",x"24",x"00",
x"00",x"42",x"24",x"18",x"18",x"24",x"42",x"00",x"00",x"82",x"44",x"28",x"10",x"10",x"10",x"00",
x"00",x"7E",x"04",x"08",x"10",x"20",x"7E",x"00",x"00",x"0E",x"08",x"08",x"08",x"08",x"0E",x"00",
x"00",x"00",x"40",x"20",x"10",x"08",x"04",x"00",x"00",x"70",x"10",x"10",x"10",x"10",x"70",x"00",
x"00",x"10",x"38",x"54",x"10",x"10",x"10",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"FF",
x"00",x"1C",x"22",x"78",x"20",x"20",x"7E",x"00",x"00",x"00",x"38",x"04",x"3C",x"44",x"3C",x"00",
x"00",x"20",x"20",x"3C",x"22",x"22",x"3C",x"00",x"00",x"00",x"1C",x"20",x"20",x"20",x"1C",x"00",
x"00",x"04",x"04",x"3C",x"44",x"44",x"3C",x"00",x"00",x"00",x"38",x"44",x"78",x"40",x"3C",x"00",
x"00",x"0C",x"10",x"18",x"10",x"10",x"10",x"00",x"00",x"00",x"3C",x"44",x"44",x"3C",x"04",x"38",
x"00",x"40",x"40",x"78",x"44",x"44",x"44",x"00",x"00",x"10",x"00",x"30",x"10",x"10",x"38",x"00",
x"00",x"04",x"00",x"04",x"04",x"04",x"24",x"18",x"00",x"20",x"28",x"30",x"30",x"28",x"24",x"00",
x"00",x"10",x"10",x"10",x"10",x"10",x"0C",x"00",x"00",x"00",x"68",x"54",x"54",x"54",x"54",x"00",
x"00",x"00",x"78",x"44",x"44",x"44",x"44",x"00",x"00",x"00",x"38",x"44",x"44",x"44",x"38",x"00",
x"00",x"00",x"78",x"44",x"44",x"78",x"40",x"40",x"00",x"00",x"3C",x"44",x"44",x"3C",x"04",x"06",
x"00",x"00",x"1C",x"20",x"20",x"20",x"20",x"00",x"00",x"00",x"38",x"40",x"38",x"04",x"78",x"00",
x"00",x"10",x"38",x"10",x"10",x"10",x"0C",x"00",x"00",x"00",x"44",x"44",x"44",x"44",x"38",x"00",
x"00",x"00",x"44",x"44",x"28",x"28",x"10",x"00",x"00",x"00",x"44",x"54",x"54",x"54",x"28",x"00",
x"00",x"00",x"44",x"28",x"10",x"28",x"44",x"00",x"00",x"00",x"44",x"44",x"44",x"3C",x"04",x"38",
x"00",x"00",x"7C",x"08",x"10",x"20",x"7C",x"00",x"00",x"0E",x"08",x"30",x"08",x"08",x"0E",x"00",
x"00",x"08",x"08",x"08",x"08",x"08",x"08",x"00",x"00",x"70",x"10",x"0C",x"10",x"10",x"70",x"00",
x"00",x"14",x"28",x"00",x"00",x"00",x"00",x"00",x"3C",x"42",x"99",x"A1",x"A1",x"99",x"42",x"3C"

);

begin

  process(CLK)
  begin
    if rising_edge(CLK) then
	   if WR='1' then
		  myROM(conv_integer(A)) <= DIN;
		end if;
	   DOUT <= myROM(conv_integer(A));
	 end if;
  end process;
  
end Behavioral;

